`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module Memo(
  input         clock,
  input         io_wen,
  input  [7:0]  io_wrAddr,
  input  [17:0] io_wrData,
  input         io_ren,
  input  [7:0]  io_rdAddr,
  output [17:0] io_rdData
);
  reg [17:0] mem [0:255];
  reg [31:0] _GEN_0;
  wire [17:0] mem__T_12_data;
  wire [7:0] mem__T_12_addr;
  wire [17:0] mem__T_10_data;
  wire [7:0] mem__T_10_addr;
  wire  mem__T_10_mask;
  wire  mem__T_10_en;
  wire [17:0] _GEN_7;
  assign io_rdData = _GEN_7;
  assign mem__T_12_addr = io_rdAddr;
  assign mem__T_12_data = mem[mem__T_12_addr];
  assign mem__T_10_data = io_wrData;
  assign mem__T_10_addr = io_wrAddr;
  assign mem__T_10_mask = io_wen;
  assign mem__T_10_en = io_wen;
  assign _GEN_7 = io_ren ? mem__T_12_data : 18'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    mem[initvar] = _GEN_0[17:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if(mem__T_10_en & mem__T_10_mask) begin
      mem[mem__T_10_addr] <= mem__T_10_data;
    end
  end
endmodule
module AggregateMem(
  input          clock,
  input  [7:0]   io_addr,
  input  [127:0] io_in,
  output [127:0] io_out,
  input          io_wen,
  input          io_ren
);
  wire  Memo_clock;
  wire  Memo_io_wen;
  wire [7:0] Memo_io_wrAddr;
  wire [17:0] Memo_io_wrData;
  wire  Memo_io_ren;
  wire [7:0] Memo_io_rdAddr;
  wire [17:0] Memo_io_rdData;
  wire  Memo_1_clock;
  wire  Memo_1_io_wen;
  wire [7:0] Memo_1_io_wrAddr;
  wire [17:0] Memo_1_io_wrData;
  wire  Memo_1_io_ren;
  wire [7:0] Memo_1_io_rdAddr;
  wire [17:0] Memo_1_io_rdData;
  wire  Memo_2_clock;
  wire  Memo_2_io_wen;
  wire [7:0] Memo_2_io_wrAddr;
  wire [17:0] Memo_2_io_wrData;
  wire  Memo_2_io_ren;
  wire [7:0] Memo_2_io_rdAddr;
  wire [17:0] Memo_2_io_rdData;
  wire  Memo_3_clock;
  wire  Memo_3_io_wen;
  wire [7:0] Memo_3_io_wrAddr;
  wire [17:0] Memo_3_io_wrData;
  wire  Memo_3_io_ren;
  wire [7:0] Memo_3_io_rdAddr;
  wire [17:0] Memo_3_io_rdData;
  wire  Memo_4_clock;
  wire  Memo_4_io_wen;
  wire [7:0] Memo_4_io_wrAddr;
  wire [17:0] Memo_4_io_wrData;
  wire  Memo_4_io_ren;
  wire [7:0] Memo_4_io_rdAddr;
  wire [17:0] Memo_4_io_rdData;
  wire  Memo_5_clock;
  wire  Memo_5_io_wen;
  wire [7:0] Memo_5_io_wrAddr;
  wire [17:0] Memo_5_io_wrData;
  wire  Memo_5_io_ren;
  wire [7:0] Memo_5_io_rdAddr;
  wire [17:0] Memo_5_io_rdData;
  wire  Memo_6_clock;
  wire  Memo_6_io_wen;
  wire [7:0] Memo_6_io_wrAddr;
  wire [17:0] Memo_6_io_wrData;
  wire  Memo_6_io_ren;
  wire [7:0] Memo_6_io_rdAddr;
  wire [17:0] Memo_6_io_rdData;
  wire  Memo_7_clock;
  wire  Memo_7_io_wen;
  wire [7:0] Memo_7_io_wrAddr;
  wire [17:0] Memo_7_io_wrData;
  wire  Memo_7_io_ren;
  wire [7:0] Memo_7_io_rdAddr;
  wire [17:0] Memo_7_io_rdData;
  wire [15:0] _T_8;
  wire [17:0] _T_9;
  wire [15:0] _T_11;
  wire [17:0] _T_12;
  wire [15:0] _T_14;
  wire [17:0] _T_15;
  wire [15:0] _T_17;
  wire [17:0] _T_18;
  wire [15:0] _T_20;
  wire [17:0] _T_21;
  wire [15:0] _T_23;
  wire [17:0] _T_24;
  wire [15:0] _T_26;
  wire [17:0] _T_27;
  wire [15:0] _T_29;
  wire [17:0] _T_30;
  wire [15:0] _T_31;
  wire [15:0] _T_32;
  wire [15:0] _T_33;
  wire [15:0] _T_34;
  wire [15:0] _T_35;
  wire [15:0] _T_36;
  wire [15:0] _T_37;
  wire [15:0] _T_38;
  wire [31:0] _T_39;
  wire [31:0] _T_40;
  wire [63:0] _T_41;
  wire [31:0] _T_42;
  wire [31:0] _T_43;
  wire [63:0] _T_44;
  wire [127:0] _T_45;
  Memo Memo (
    .clock(Memo_clock),
    .io_wen(Memo_io_wen),
    .io_wrAddr(Memo_io_wrAddr),
    .io_wrData(Memo_io_wrData),
    .io_ren(Memo_io_ren),
    .io_rdAddr(Memo_io_rdAddr),
    .io_rdData(Memo_io_rdData)
  );
  Memo Memo_1 (
    .clock(Memo_1_clock),
    .io_wen(Memo_1_io_wen),
    .io_wrAddr(Memo_1_io_wrAddr),
    .io_wrData(Memo_1_io_wrData),
    .io_ren(Memo_1_io_ren),
    .io_rdAddr(Memo_1_io_rdAddr),
    .io_rdData(Memo_1_io_rdData)
  );
  Memo Memo_2 (
    .clock(Memo_2_clock),
    .io_wen(Memo_2_io_wen),
    .io_wrAddr(Memo_2_io_wrAddr),
    .io_wrData(Memo_2_io_wrData),
    .io_ren(Memo_2_io_ren),
    .io_rdAddr(Memo_2_io_rdAddr),
    .io_rdData(Memo_2_io_rdData)
  );
  Memo Memo_3 (
    .clock(Memo_3_clock),
    .io_wen(Memo_3_io_wen),
    .io_wrAddr(Memo_3_io_wrAddr),
    .io_wrData(Memo_3_io_wrData),
    .io_ren(Memo_3_io_ren),
    .io_rdAddr(Memo_3_io_rdAddr),
    .io_rdData(Memo_3_io_rdData)
  );
  Memo Memo_4 (
    .clock(Memo_4_clock),
    .io_wen(Memo_4_io_wen),
    .io_wrAddr(Memo_4_io_wrAddr),
    .io_wrData(Memo_4_io_wrData),
    .io_ren(Memo_4_io_ren),
    .io_rdAddr(Memo_4_io_rdAddr),
    .io_rdData(Memo_4_io_rdData)
  );
  Memo Memo_5 (
    .clock(Memo_5_clock),
    .io_wen(Memo_5_io_wen),
    .io_wrAddr(Memo_5_io_wrAddr),
    .io_wrData(Memo_5_io_wrData),
    .io_ren(Memo_5_io_ren),
    .io_rdAddr(Memo_5_io_rdAddr),
    .io_rdData(Memo_5_io_rdData)
  );
  Memo Memo_6 (
    .clock(Memo_6_clock),
    .io_wen(Memo_6_io_wen),
    .io_wrAddr(Memo_6_io_wrAddr),
    .io_wrData(Memo_6_io_wrData),
    .io_ren(Memo_6_io_ren),
    .io_rdAddr(Memo_6_io_rdAddr),
    .io_rdData(Memo_6_io_rdData)
  );
  Memo Memo_7 (
    .clock(Memo_7_clock),
    .io_wen(Memo_7_io_wen),
    .io_wrAddr(Memo_7_io_wrAddr),
    .io_wrData(Memo_7_io_wrData),
    .io_ren(Memo_7_io_ren),
    .io_rdAddr(Memo_7_io_rdAddr),
    .io_rdData(Memo_7_io_rdData)
  );
  assign io_out = _T_45;
  assign Memo_clock = clock;
  assign Memo_io_wen = io_wen;
  assign Memo_io_wrAddr = io_addr;
  assign Memo_io_wrData = _T_9;
  assign Memo_io_ren = io_ren;
  assign Memo_io_rdAddr = io_addr;
  assign Memo_1_clock = clock;
  assign Memo_1_io_wen = io_wen;
  assign Memo_1_io_wrAddr = io_addr;
  assign Memo_1_io_wrData = _T_12;
  assign Memo_1_io_ren = io_ren;
  assign Memo_1_io_rdAddr = io_addr;
  assign Memo_2_clock = clock;
  assign Memo_2_io_wen = io_wen;
  assign Memo_2_io_wrAddr = io_addr;
  assign Memo_2_io_wrData = _T_15;
  assign Memo_2_io_ren = io_ren;
  assign Memo_2_io_rdAddr = io_addr;
  assign Memo_3_clock = clock;
  assign Memo_3_io_wen = io_wen;
  assign Memo_3_io_wrAddr = io_addr;
  assign Memo_3_io_wrData = _T_18;
  assign Memo_3_io_ren = io_ren;
  assign Memo_3_io_rdAddr = io_addr;
  assign Memo_4_clock = clock;
  assign Memo_4_io_wen = io_wen;
  assign Memo_4_io_wrAddr = io_addr;
  assign Memo_4_io_wrData = _T_21;
  assign Memo_4_io_ren = io_ren;
  assign Memo_4_io_rdAddr = io_addr;
  assign Memo_5_clock = clock;
  assign Memo_5_io_wen = io_wen;
  assign Memo_5_io_wrAddr = io_addr;
  assign Memo_5_io_wrData = _T_24;
  assign Memo_5_io_ren = io_ren;
  assign Memo_5_io_rdAddr = io_addr;
  assign Memo_6_clock = clock;
  assign Memo_6_io_wen = io_wen;
  assign Memo_6_io_wrAddr = io_addr;
  assign Memo_6_io_wrData = _T_27;
  assign Memo_6_io_ren = io_ren;
  assign Memo_6_io_rdAddr = io_addr;
  assign Memo_7_clock = clock;
  assign Memo_7_io_wen = io_wen;
  assign Memo_7_io_wrAddr = io_addr;
  assign Memo_7_io_wrData = _T_30;
  assign Memo_7_io_ren = io_ren;
  assign Memo_7_io_rdAddr = io_addr;
  assign _T_8 = io_in[15:0];
  assign _T_9 = {2'h0,_T_8};
  assign _T_11 = io_in[31:16];
  assign _T_12 = {2'h0,_T_11};
  assign _T_14 = io_in[47:32];
  assign _T_15 = {2'h0,_T_14};
  assign _T_17 = io_in[63:48];
  assign _T_18 = {2'h0,_T_17};
  assign _T_20 = io_in[79:64];
  assign _T_21 = {2'h0,_T_20};
  assign _T_23 = io_in[95:80];
  assign _T_24 = {2'h0,_T_23};
  assign _T_26 = io_in[111:96];
  assign _T_27 = {2'h0,_T_26};
  assign _T_29 = io_in[127:112];
  assign _T_30 = {2'h0,_T_29};
  assign _T_31 = Memo_7_io_rdData[15:0];
  assign _T_32 = Memo_6_io_rdData[15:0];
  assign _T_33 = Memo_5_io_rdData[15:0];
  assign _T_34 = Memo_4_io_rdData[15:0];
  assign _T_35 = Memo_3_io_rdData[15:0];
  assign _T_36 = Memo_2_io_rdData[15:0];
  assign _T_37 = Memo_1_io_rdData[15:0];
  assign _T_38 = Memo_io_rdData[15:0];
  assign _T_39 = {_T_37,_T_38};
  assign _T_40 = {_T_35,_T_36};
  assign _T_41 = {_T_40,_T_39};
  assign _T_42 = {_T_33,_T_34};
  assign _T_43 = {_T_31,_T_32};
  assign _T_44 = {_T_43,_T_42};
  assign _T_45 = {_T_44,_T_41};
endmodule
module BinaryBuffer(
  input         clock,
  input         reset,
  input  [3:0]  io_in,
  input         io_push,
  output [31:0] io_out,
  input         io_pop
);
  reg [5:0] wPos;
  reg [31:0] _GEN_139;
  reg [2:0] rPos;
  reg [31:0] _GEN_140;
  reg [3:0] mem_0;
  reg [31:0] _GEN_141;
  reg [3:0] mem_1;
  reg [31:0] _GEN_142;
  reg [3:0] mem_2;
  reg [31:0] _GEN_143;
  reg [3:0] mem_3;
  reg [31:0] _GEN_144;
  reg [3:0] mem_4;
  reg [31:0] _GEN_145;
  reg [3:0] mem_5;
  reg [31:0] _GEN_146;
  reg [3:0] mem_6;
  reg [31:0] _GEN_147;
  reg [3:0] mem_7;
  reg [31:0] _GEN_148;
  reg [3:0] mem_8;
  reg [31:0] _GEN_149;
  reg [3:0] mem_9;
  reg [31:0] _GEN_150;
  reg [3:0] mem_10;
  reg [31:0] _GEN_151;
  reg [3:0] mem_11;
  reg [31:0] _GEN_152;
  reg [3:0] mem_12;
  reg [31:0] _GEN_153;
  reg [3:0] mem_13;
  reg [31:0] _GEN_154;
  reg [3:0] mem_14;
  reg [31:0] _GEN_155;
  reg [3:0] mem_15;
  reg [31:0] _GEN_156;
  reg [3:0] mem_16;
  reg [31:0] _GEN_157;
  reg [3:0] mem_17;
  reg [31:0] _GEN_158;
  reg [3:0] mem_18;
  reg [31:0] _GEN_159;
  reg [3:0] mem_19;
  reg [31:0] _GEN_160;
  reg [3:0] mem_20;
  reg [31:0] _GEN_161;
  reg [3:0] mem_21;
  reg [31:0] _GEN_162;
  reg [3:0] mem_22;
  reg [31:0] _GEN_163;
  reg [3:0] mem_23;
  reg [31:0] _GEN_164;
  reg [3:0] mem_24;
  reg [31:0] _GEN_165;
  reg [3:0] mem_25;
  reg [31:0] _GEN_166;
  reg [3:0] mem_26;
  reg [31:0] _GEN_167;
  reg [3:0] mem_27;
  reg [31:0] _GEN_168;
  reg [3:0] mem_28;
  reg [31:0] _GEN_169;
  reg [3:0] mem_29;
  reg [31:0] _GEN_170;
  reg [3:0] mem_30;
  reg [31:0] _GEN_171;
  reg [3:0] mem_31;
  reg [31:0] _GEN_172;
  reg [3:0] mem_32;
  reg [31:0] _GEN_173;
  reg [3:0] mem_33;
  reg [31:0] _GEN_174;
  reg [3:0] mem_34;
  reg [31:0] _GEN_175;
  reg [3:0] mem_35;
  reg [31:0] _GEN_176;
  reg [3:0] mem_36;
  reg [31:0] _GEN_177;
  reg [3:0] mem_37;
  reg [31:0] _GEN_178;
  reg [3:0] mem_38;
  reg [31:0] _GEN_179;
  reg [3:0] mem_39;
  reg [31:0] _GEN_180;
  reg [3:0] mem_40;
  reg [31:0] _GEN_181;
  reg [3:0] mem_41;
  reg [31:0] _GEN_182;
  reg [3:0] mem_42;
  reg [31:0] _GEN_183;
  reg [3:0] mem_43;
  reg [31:0] _GEN_184;
  reg [3:0] mem_44;
  reg [31:0] _GEN_185;
  reg [3:0] mem_45;
  reg [31:0] _GEN_186;
  reg [3:0] mem_46;
  reg [31:0] _GEN_187;
  reg [3:0] mem_47;
  reg [31:0] _GEN_188;
  reg [3:0] mem_48;
  reg [31:0] _GEN_189;
  reg [3:0] mem_49;
  reg [31:0] _GEN_190;
  reg [3:0] mem_50;
  reg [31:0] _GEN_191;
  reg [3:0] mem_51;
  reg [31:0] _GEN_192;
  reg [3:0] mem_52;
  reg [31:0] _GEN_193;
  reg [3:0] mem_53;
  reg [31:0] _GEN_194;
  reg [3:0] mem_54;
  reg [31:0] _GEN_195;
  reg [3:0] mem_55;
  reg [31:0] _GEN_196;
  reg [3:0] mem_56;
  reg [31:0] _GEN_197;
  reg [3:0] mem_57;
  reg [31:0] _GEN_198;
  reg [3:0] mem_58;
  reg [31:0] _GEN_199;
  reg [3:0] mem_59;
  reg [31:0] _GEN_200;
  reg [3:0] mem_60;
  reg [31:0] _GEN_201;
  reg [3:0] mem_61;
  reg [31:0] _GEN_202;
  reg [3:0] mem_62;
  reg [31:0] _GEN_203;
  reg [3:0] mem_63;
  reg [31:0] _GEN_204;
  wire [7:0] _T_79;
  wire [7:0] _T_80;
  wire [15:0] _T_81;
  wire [7:0] _T_82;
  wire [7:0] _T_83;
  wire [15:0] _T_84;
  wire [31:0] _T_85;
  wire [7:0] _T_86;
  wire [7:0] _T_87;
  wire [15:0] _T_88;
  wire [7:0] _T_89;
  wire [7:0] _T_90;
  wire [15:0] _T_91;
  wire [31:0] _T_92;
  wire [7:0] _T_93;
  wire [7:0] _T_94;
  wire [15:0] _T_95;
  wire [7:0] _T_96;
  wire [7:0] _T_97;
  wire [15:0] _T_98;
  wire [31:0] _T_99;
  wire [7:0] _T_100;
  wire [7:0] _T_101;
  wire [15:0] _T_102;
  wire [7:0] _T_103;
  wire [7:0] _T_104;
  wire [15:0] _T_105;
  wire [31:0] _T_106;
  wire [7:0] _T_107;
  wire [7:0] _T_108;
  wire [15:0] _T_109;
  wire [7:0] _T_110;
  wire [7:0] _T_111;
  wire [15:0] _T_112;
  wire [31:0] _T_113;
  wire [7:0] _T_114;
  wire [7:0] _T_115;
  wire [15:0] _T_116;
  wire [7:0] _T_117;
  wire [7:0] _T_118;
  wire [15:0] _T_119;
  wire [31:0] _T_120;
  wire [7:0] _T_121;
  wire [7:0] _T_122;
  wire [15:0] _T_123;
  wire [7:0] _T_124;
  wire [7:0] _T_125;
  wire [15:0] _T_126;
  wire [31:0] _T_127;
  wire [7:0] _T_128;
  wire [7:0] _T_129;
  wire [15:0] _T_130;
  wire [7:0] _T_131;
  wire [7:0] _T_132;
  wire [15:0] _T_133;
  wire [31:0] _T_134;
  wire [31:0] catMem_0;
  wire [31:0] catMem_1;
  wire [31:0] catMem_2;
  wire [31:0] catMem_3;
  wire [31:0] catMem_4;
  wire [31:0] catMem_5;
  wire [31:0] catMem_6;
  wire [31:0] catMem_7;
  wire [3:0] _GEN_0;
  wire [3:0] _GEN_2;
  wire [3:0] _GEN_3;
  wire [3:0] _GEN_4;
  wire [3:0] _GEN_5;
  wire [3:0] _GEN_6;
  wire [3:0] _GEN_7;
  wire [3:0] _GEN_8;
  wire [3:0] _GEN_9;
  wire [3:0] _GEN_10;
  wire [3:0] _GEN_11;
  wire [3:0] _GEN_12;
  wire [3:0] _GEN_13;
  wire [3:0] _GEN_14;
  wire [3:0] _GEN_15;
  wire [3:0] _GEN_16;
  wire [3:0] _GEN_17;
  wire [3:0] _GEN_18;
  wire [3:0] _GEN_19;
  wire [3:0] _GEN_20;
  wire [3:0] _GEN_21;
  wire [3:0] _GEN_22;
  wire [3:0] _GEN_23;
  wire [3:0] _GEN_24;
  wire [3:0] _GEN_25;
  wire [3:0] _GEN_26;
  wire [3:0] _GEN_27;
  wire [3:0] _GEN_28;
  wire [3:0] _GEN_29;
  wire [3:0] _GEN_30;
  wire [3:0] _GEN_31;
  wire [3:0] _GEN_32;
  wire [3:0] _GEN_33;
  wire [3:0] _GEN_34;
  wire [3:0] _GEN_35;
  wire [3:0] _GEN_36;
  wire [3:0] _GEN_37;
  wire [3:0] _GEN_38;
  wire [3:0] _GEN_39;
  wire [3:0] _GEN_40;
  wire [3:0] _GEN_41;
  wire [3:0] _GEN_42;
  wire [3:0] _GEN_43;
  wire [3:0] _GEN_44;
  wire [3:0] _GEN_45;
  wire [3:0] _GEN_46;
  wire [3:0] _GEN_47;
  wire [3:0] _GEN_48;
  wire [3:0] _GEN_49;
  wire [3:0] _GEN_50;
  wire [3:0] _GEN_51;
  wire [3:0] _GEN_52;
  wire [3:0] _GEN_53;
  wire [3:0] _GEN_54;
  wire [3:0] _GEN_55;
  wire [3:0] _GEN_56;
  wire [3:0] _GEN_57;
  wire [3:0] _GEN_58;
  wire [3:0] _GEN_59;
  wire [3:0] _GEN_60;
  wire [3:0] _GEN_61;
  wire [3:0] _GEN_62;
  wire [3:0] _GEN_63;
  wire [3:0] _GEN_64;
  wire [3:0] _GEN_65;
  wire [6:0] _T_149;
  wire [5:0] _T_150;
  wire [3:0] _GEN_66;
  wire [3:0] _GEN_67;
  wire [3:0] _GEN_68;
  wire [3:0] _GEN_69;
  wire [3:0] _GEN_70;
  wire [3:0] _GEN_71;
  wire [3:0] _GEN_72;
  wire [3:0] _GEN_73;
  wire [3:0] _GEN_74;
  wire [3:0] _GEN_75;
  wire [3:0] _GEN_76;
  wire [3:0] _GEN_77;
  wire [3:0] _GEN_78;
  wire [3:0] _GEN_79;
  wire [3:0] _GEN_80;
  wire [3:0] _GEN_81;
  wire [3:0] _GEN_82;
  wire [3:0] _GEN_83;
  wire [3:0] _GEN_84;
  wire [3:0] _GEN_85;
  wire [3:0] _GEN_86;
  wire [3:0] _GEN_87;
  wire [3:0] _GEN_88;
  wire [3:0] _GEN_89;
  wire [3:0] _GEN_90;
  wire [3:0] _GEN_91;
  wire [3:0] _GEN_92;
  wire [3:0] _GEN_93;
  wire [3:0] _GEN_94;
  wire [3:0] _GEN_95;
  wire [3:0] _GEN_96;
  wire [3:0] _GEN_97;
  wire [3:0] _GEN_98;
  wire [3:0] _GEN_99;
  wire [3:0] _GEN_100;
  wire [3:0] _GEN_101;
  wire [3:0] _GEN_102;
  wire [3:0] _GEN_103;
  wire [3:0] _GEN_104;
  wire [3:0] _GEN_105;
  wire [3:0] _GEN_106;
  wire [3:0] _GEN_107;
  wire [3:0] _GEN_108;
  wire [3:0] _GEN_109;
  wire [3:0] _GEN_110;
  wire [3:0] _GEN_111;
  wire [3:0] _GEN_112;
  wire [3:0] _GEN_113;
  wire [3:0] _GEN_114;
  wire [3:0] _GEN_115;
  wire [3:0] _GEN_116;
  wire [3:0] _GEN_117;
  wire [3:0] _GEN_118;
  wire [3:0] _GEN_119;
  wire [3:0] _GEN_120;
  wire [3:0] _GEN_121;
  wire [3:0] _GEN_122;
  wire [3:0] _GEN_123;
  wire [3:0] _GEN_124;
  wire [3:0] _GEN_125;
  wire [3:0] _GEN_126;
  wire [3:0] _GEN_127;
  wire [3:0] _GEN_128;
  wire [3:0] _GEN_129;
  wire [5:0] _GEN_130;
  wire [3:0] _T_152;
  wire [2:0] _T_153;
  wire [2:0] _GEN_131;
  wire [31:0] _GEN_1;
  wire [31:0] _GEN_132;
  wire [31:0] _GEN_133;
  wire [31:0] _GEN_134;
  wire [31:0] _GEN_135;
  wire [31:0] _GEN_136;
  wire [31:0] _GEN_137;
  wire [31:0] _GEN_138;
  assign io_out = _GEN_1;
  assign _T_79 = {mem_6,mem_7};
  assign _T_80 = {mem_4,mem_5};
  assign _T_81 = {_T_80,_T_79};
  assign _T_82 = {mem_2,mem_3};
  assign _T_83 = {mem_0,mem_1};
  assign _T_84 = {_T_83,_T_82};
  assign _T_85 = {_T_84,_T_81};
  assign _T_86 = {mem_14,mem_15};
  assign _T_87 = {mem_12,mem_13};
  assign _T_88 = {_T_87,_T_86};
  assign _T_89 = {mem_10,mem_11};
  assign _T_90 = {mem_8,mem_9};
  assign _T_91 = {_T_90,_T_89};
  assign _T_92 = {_T_91,_T_88};
  assign _T_93 = {mem_22,mem_23};
  assign _T_94 = {mem_20,mem_21};
  assign _T_95 = {_T_94,_T_93};
  assign _T_96 = {mem_18,mem_19};
  assign _T_97 = {mem_16,mem_17};
  assign _T_98 = {_T_97,_T_96};
  assign _T_99 = {_T_98,_T_95};
  assign _T_100 = {mem_30,mem_31};
  assign _T_101 = {mem_28,mem_29};
  assign _T_102 = {_T_101,_T_100};
  assign _T_103 = {mem_26,mem_27};
  assign _T_104 = {mem_24,mem_25};
  assign _T_105 = {_T_104,_T_103};
  assign _T_106 = {_T_105,_T_102};
  assign _T_107 = {mem_38,mem_39};
  assign _T_108 = {mem_36,mem_37};
  assign _T_109 = {_T_108,_T_107};
  assign _T_110 = {mem_34,mem_35};
  assign _T_111 = {mem_32,mem_33};
  assign _T_112 = {_T_111,_T_110};
  assign _T_113 = {_T_112,_T_109};
  assign _T_114 = {mem_46,mem_47};
  assign _T_115 = {mem_44,mem_45};
  assign _T_116 = {_T_115,_T_114};
  assign _T_117 = {mem_42,mem_43};
  assign _T_118 = {mem_40,mem_41};
  assign _T_119 = {_T_118,_T_117};
  assign _T_120 = {_T_119,_T_116};
  assign _T_121 = {mem_54,mem_55};
  assign _T_122 = {mem_52,mem_53};
  assign _T_123 = {_T_122,_T_121};
  assign _T_124 = {mem_50,mem_51};
  assign _T_125 = {mem_48,mem_49};
  assign _T_126 = {_T_125,_T_124};
  assign _T_127 = {_T_126,_T_123};
  assign _T_128 = {mem_62,mem_63};
  assign _T_129 = {mem_60,mem_61};
  assign _T_130 = {_T_129,_T_128};
  assign _T_131 = {mem_58,mem_59};
  assign _T_132 = {mem_56,mem_57};
  assign _T_133 = {_T_132,_T_131};
  assign _T_134 = {_T_133,_T_130};
  assign catMem_0 = _T_85;
  assign catMem_1 = _T_92;
  assign catMem_2 = _T_99;
  assign catMem_3 = _T_106;
  assign catMem_4 = _T_113;
  assign catMem_5 = _T_120;
  assign catMem_6 = _T_127;
  assign catMem_7 = _T_134;
  assign _GEN_0 = io_in;
  assign _GEN_2 = 6'h0 == wPos ? _GEN_0 : mem_0;
  assign _GEN_3 = 6'h1 == wPos ? _GEN_0 : mem_1;
  assign _GEN_4 = 6'h2 == wPos ? _GEN_0 : mem_2;
  assign _GEN_5 = 6'h3 == wPos ? _GEN_0 : mem_3;
  assign _GEN_6 = 6'h4 == wPos ? _GEN_0 : mem_4;
  assign _GEN_7 = 6'h5 == wPos ? _GEN_0 : mem_5;
  assign _GEN_8 = 6'h6 == wPos ? _GEN_0 : mem_6;
  assign _GEN_9 = 6'h7 == wPos ? _GEN_0 : mem_7;
  assign _GEN_10 = 6'h8 == wPos ? _GEN_0 : mem_8;
  assign _GEN_11 = 6'h9 == wPos ? _GEN_0 : mem_9;
  assign _GEN_12 = 6'ha == wPos ? _GEN_0 : mem_10;
  assign _GEN_13 = 6'hb == wPos ? _GEN_0 : mem_11;
  assign _GEN_14 = 6'hc == wPos ? _GEN_0 : mem_12;
  assign _GEN_15 = 6'hd == wPos ? _GEN_0 : mem_13;
  assign _GEN_16 = 6'he == wPos ? _GEN_0 : mem_14;
  assign _GEN_17 = 6'hf == wPos ? _GEN_0 : mem_15;
  assign _GEN_18 = 6'h10 == wPos ? _GEN_0 : mem_16;
  assign _GEN_19 = 6'h11 == wPos ? _GEN_0 : mem_17;
  assign _GEN_20 = 6'h12 == wPos ? _GEN_0 : mem_18;
  assign _GEN_21 = 6'h13 == wPos ? _GEN_0 : mem_19;
  assign _GEN_22 = 6'h14 == wPos ? _GEN_0 : mem_20;
  assign _GEN_23 = 6'h15 == wPos ? _GEN_0 : mem_21;
  assign _GEN_24 = 6'h16 == wPos ? _GEN_0 : mem_22;
  assign _GEN_25 = 6'h17 == wPos ? _GEN_0 : mem_23;
  assign _GEN_26 = 6'h18 == wPos ? _GEN_0 : mem_24;
  assign _GEN_27 = 6'h19 == wPos ? _GEN_0 : mem_25;
  assign _GEN_28 = 6'h1a == wPos ? _GEN_0 : mem_26;
  assign _GEN_29 = 6'h1b == wPos ? _GEN_0 : mem_27;
  assign _GEN_30 = 6'h1c == wPos ? _GEN_0 : mem_28;
  assign _GEN_31 = 6'h1d == wPos ? _GEN_0 : mem_29;
  assign _GEN_32 = 6'h1e == wPos ? _GEN_0 : mem_30;
  assign _GEN_33 = 6'h1f == wPos ? _GEN_0 : mem_31;
  assign _GEN_34 = 6'h20 == wPos ? _GEN_0 : mem_32;
  assign _GEN_35 = 6'h21 == wPos ? _GEN_0 : mem_33;
  assign _GEN_36 = 6'h22 == wPos ? _GEN_0 : mem_34;
  assign _GEN_37 = 6'h23 == wPos ? _GEN_0 : mem_35;
  assign _GEN_38 = 6'h24 == wPos ? _GEN_0 : mem_36;
  assign _GEN_39 = 6'h25 == wPos ? _GEN_0 : mem_37;
  assign _GEN_40 = 6'h26 == wPos ? _GEN_0 : mem_38;
  assign _GEN_41 = 6'h27 == wPos ? _GEN_0 : mem_39;
  assign _GEN_42 = 6'h28 == wPos ? _GEN_0 : mem_40;
  assign _GEN_43 = 6'h29 == wPos ? _GEN_0 : mem_41;
  assign _GEN_44 = 6'h2a == wPos ? _GEN_0 : mem_42;
  assign _GEN_45 = 6'h2b == wPos ? _GEN_0 : mem_43;
  assign _GEN_46 = 6'h2c == wPos ? _GEN_0 : mem_44;
  assign _GEN_47 = 6'h2d == wPos ? _GEN_0 : mem_45;
  assign _GEN_48 = 6'h2e == wPos ? _GEN_0 : mem_46;
  assign _GEN_49 = 6'h2f == wPos ? _GEN_0 : mem_47;
  assign _GEN_50 = 6'h30 == wPos ? _GEN_0 : mem_48;
  assign _GEN_51 = 6'h31 == wPos ? _GEN_0 : mem_49;
  assign _GEN_52 = 6'h32 == wPos ? _GEN_0 : mem_50;
  assign _GEN_53 = 6'h33 == wPos ? _GEN_0 : mem_51;
  assign _GEN_54 = 6'h34 == wPos ? _GEN_0 : mem_52;
  assign _GEN_55 = 6'h35 == wPos ? _GEN_0 : mem_53;
  assign _GEN_56 = 6'h36 == wPos ? _GEN_0 : mem_54;
  assign _GEN_57 = 6'h37 == wPos ? _GEN_0 : mem_55;
  assign _GEN_58 = 6'h38 == wPos ? _GEN_0 : mem_56;
  assign _GEN_59 = 6'h39 == wPos ? _GEN_0 : mem_57;
  assign _GEN_60 = 6'h3a == wPos ? _GEN_0 : mem_58;
  assign _GEN_61 = 6'h3b == wPos ? _GEN_0 : mem_59;
  assign _GEN_62 = 6'h3c == wPos ? _GEN_0 : mem_60;
  assign _GEN_63 = 6'h3d == wPos ? _GEN_0 : mem_61;
  assign _GEN_64 = 6'h3e == wPos ? _GEN_0 : mem_62;
  assign _GEN_65 = 6'h3f == wPos ? _GEN_0 : mem_63;
  assign _T_149 = wPos + 6'h1;
  assign _T_150 = _T_149[5:0];
  assign _GEN_66 = io_push ? _GEN_2 : mem_0;
  assign _GEN_67 = io_push ? _GEN_3 : mem_1;
  assign _GEN_68 = io_push ? _GEN_4 : mem_2;
  assign _GEN_69 = io_push ? _GEN_5 : mem_3;
  assign _GEN_70 = io_push ? _GEN_6 : mem_4;
  assign _GEN_71 = io_push ? _GEN_7 : mem_5;
  assign _GEN_72 = io_push ? _GEN_8 : mem_6;
  assign _GEN_73 = io_push ? _GEN_9 : mem_7;
  assign _GEN_74 = io_push ? _GEN_10 : mem_8;
  assign _GEN_75 = io_push ? _GEN_11 : mem_9;
  assign _GEN_76 = io_push ? _GEN_12 : mem_10;
  assign _GEN_77 = io_push ? _GEN_13 : mem_11;
  assign _GEN_78 = io_push ? _GEN_14 : mem_12;
  assign _GEN_79 = io_push ? _GEN_15 : mem_13;
  assign _GEN_80 = io_push ? _GEN_16 : mem_14;
  assign _GEN_81 = io_push ? _GEN_17 : mem_15;
  assign _GEN_82 = io_push ? _GEN_18 : mem_16;
  assign _GEN_83 = io_push ? _GEN_19 : mem_17;
  assign _GEN_84 = io_push ? _GEN_20 : mem_18;
  assign _GEN_85 = io_push ? _GEN_21 : mem_19;
  assign _GEN_86 = io_push ? _GEN_22 : mem_20;
  assign _GEN_87 = io_push ? _GEN_23 : mem_21;
  assign _GEN_88 = io_push ? _GEN_24 : mem_22;
  assign _GEN_89 = io_push ? _GEN_25 : mem_23;
  assign _GEN_90 = io_push ? _GEN_26 : mem_24;
  assign _GEN_91 = io_push ? _GEN_27 : mem_25;
  assign _GEN_92 = io_push ? _GEN_28 : mem_26;
  assign _GEN_93 = io_push ? _GEN_29 : mem_27;
  assign _GEN_94 = io_push ? _GEN_30 : mem_28;
  assign _GEN_95 = io_push ? _GEN_31 : mem_29;
  assign _GEN_96 = io_push ? _GEN_32 : mem_30;
  assign _GEN_97 = io_push ? _GEN_33 : mem_31;
  assign _GEN_98 = io_push ? _GEN_34 : mem_32;
  assign _GEN_99 = io_push ? _GEN_35 : mem_33;
  assign _GEN_100 = io_push ? _GEN_36 : mem_34;
  assign _GEN_101 = io_push ? _GEN_37 : mem_35;
  assign _GEN_102 = io_push ? _GEN_38 : mem_36;
  assign _GEN_103 = io_push ? _GEN_39 : mem_37;
  assign _GEN_104 = io_push ? _GEN_40 : mem_38;
  assign _GEN_105 = io_push ? _GEN_41 : mem_39;
  assign _GEN_106 = io_push ? _GEN_42 : mem_40;
  assign _GEN_107 = io_push ? _GEN_43 : mem_41;
  assign _GEN_108 = io_push ? _GEN_44 : mem_42;
  assign _GEN_109 = io_push ? _GEN_45 : mem_43;
  assign _GEN_110 = io_push ? _GEN_46 : mem_44;
  assign _GEN_111 = io_push ? _GEN_47 : mem_45;
  assign _GEN_112 = io_push ? _GEN_48 : mem_46;
  assign _GEN_113 = io_push ? _GEN_49 : mem_47;
  assign _GEN_114 = io_push ? _GEN_50 : mem_48;
  assign _GEN_115 = io_push ? _GEN_51 : mem_49;
  assign _GEN_116 = io_push ? _GEN_52 : mem_50;
  assign _GEN_117 = io_push ? _GEN_53 : mem_51;
  assign _GEN_118 = io_push ? _GEN_54 : mem_52;
  assign _GEN_119 = io_push ? _GEN_55 : mem_53;
  assign _GEN_120 = io_push ? _GEN_56 : mem_54;
  assign _GEN_121 = io_push ? _GEN_57 : mem_55;
  assign _GEN_122 = io_push ? _GEN_58 : mem_56;
  assign _GEN_123 = io_push ? _GEN_59 : mem_57;
  assign _GEN_124 = io_push ? _GEN_60 : mem_58;
  assign _GEN_125 = io_push ? _GEN_61 : mem_59;
  assign _GEN_126 = io_push ? _GEN_62 : mem_60;
  assign _GEN_127 = io_push ? _GEN_63 : mem_61;
  assign _GEN_128 = io_push ? _GEN_64 : mem_62;
  assign _GEN_129 = io_push ? _GEN_65 : mem_63;
  assign _GEN_130 = io_push ? _T_150 : wPos;
  assign _T_152 = rPos + 3'h1;
  assign _T_153 = _T_152[2:0];
  assign _GEN_131 = io_pop ? _T_153 : rPos;
  assign _GEN_1 = _GEN_138;
  assign _GEN_132 = 3'h1 == rPos ? catMem_1 : catMem_0;
  assign _GEN_133 = 3'h2 == rPos ? catMem_2 : _GEN_132;
  assign _GEN_134 = 3'h3 == rPos ? catMem_3 : _GEN_133;
  assign _GEN_135 = 3'h4 == rPos ? catMem_4 : _GEN_134;
  assign _GEN_136 = 3'h5 == rPos ? catMem_5 : _GEN_135;
  assign _GEN_137 = 3'h6 == rPos ? catMem_6 : _GEN_136;
  assign _GEN_138 = 3'h7 == rPos ? catMem_7 : _GEN_137;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_139 = {1{$random}};
  wPos = _GEN_139[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_140 = {1{$random}};
  rPos = _GEN_140[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_141 = {1{$random}};
  mem_0 = _GEN_141[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_142 = {1{$random}};
  mem_1 = _GEN_142[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_143 = {1{$random}};
  mem_2 = _GEN_143[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_144 = {1{$random}};
  mem_3 = _GEN_144[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_145 = {1{$random}};
  mem_4 = _GEN_145[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_146 = {1{$random}};
  mem_5 = _GEN_146[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_147 = {1{$random}};
  mem_6 = _GEN_147[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_148 = {1{$random}};
  mem_7 = _GEN_148[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_149 = {1{$random}};
  mem_8 = _GEN_149[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_150 = {1{$random}};
  mem_9 = _GEN_150[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_151 = {1{$random}};
  mem_10 = _GEN_151[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_152 = {1{$random}};
  mem_11 = _GEN_152[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_153 = {1{$random}};
  mem_12 = _GEN_153[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_154 = {1{$random}};
  mem_13 = _GEN_154[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_155 = {1{$random}};
  mem_14 = _GEN_155[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_156 = {1{$random}};
  mem_15 = _GEN_156[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_157 = {1{$random}};
  mem_16 = _GEN_157[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_158 = {1{$random}};
  mem_17 = _GEN_158[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_159 = {1{$random}};
  mem_18 = _GEN_159[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_160 = {1{$random}};
  mem_19 = _GEN_160[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_161 = {1{$random}};
  mem_20 = _GEN_161[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_162 = {1{$random}};
  mem_21 = _GEN_162[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_163 = {1{$random}};
  mem_22 = _GEN_163[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_164 = {1{$random}};
  mem_23 = _GEN_164[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_165 = {1{$random}};
  mem_24 = _GEN_165[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_166 = {1{$random}};
  mem_25 = _GEN_166[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_167 = {1{$random}};
  mem_26 = _GEN_167[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_168 = {1{$random}};
  mem_27 = _GEN_168[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_169 = {1{$random}};
  mem_28 = _GEN_169[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_170 = {1{$random}};
  mem_29 = _GEN_170[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_171 = {1{$random}};
  mem_30 = _GEN_171[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_172 = {1{$random}};
  mem_31 = _GEN_172[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_173 = {1{$random}};
  mem_32 = _GEN_173[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_174 = {1{$random}};
  mem_33 = _GEN_174[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_175 = {1{$random}};
  mem_34 = _GEN_175[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_176 = {1{$random}};
  mem_35 = _GEN_176[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_177 = {1{$random}};
  mem_36 = _GEN_177[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_178 = {1{$random}};
  mem_37 = _GEN_178[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_179 = {1{$random}};
  mem_38 = _GEN_179[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_180 = {1{$random}};
  mem_39 = _GEN_180[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_181 = {1{$random}};
  mem_40 = _GEN_181[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_182 = {1{$random}};
  mem_41 = _GEN_182[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_183 = {1{$random}};
  mem_42 = _GEN_183[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_184 = {1{$random}};
  mem_43 = _GEN_184[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_185 = {1{$random}};
  mem_44 = _GEN_185[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_186 = {1{$random}};
  mem_45 = _GEN_186[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_187 = {1{$random}};
  mem_46 = _GEN_187[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_188 = {1{$random}};
  mem_47 = _GEN_188[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_189 = {1{$random}};
  mem_48 = _GEN_189[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_190 = {1{$random}};
  mem_49 = _GEN_190[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_191 = {1{$random}};
  mem_50 = _GEN_191[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_192 = {1{$random}};
  mem_51 = _GEN_192[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_193 = {1{$random}};
  mem_52 = _GEN_193[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_194 = {1{$random}};
  mem_53 = _GEN_194[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_195 = {1{$random}};
  mem_54 = _GEN_195[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_196 = {1{$random}};
  mem_55 = _GEN_196[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_197 = {1{$random}};
  mem_56 = _GEN_197[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_198 = {1{$random}};
  mem_57 = _GEN_198[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_199 = {1{$random}};
  mem_58 = _GEN_199[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_200 = {1{$random}};
  mem_59 = _GEN_200[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_201 = {1{$random}};
  mem_60 = _GEN_201[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_202 = {1{$random}};
  mem_61 = _GEN_202[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_203 = {1{$random}};
  mem_62 = _GEN_203[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_204 = {1{$random}};
  mem_63 = _GEN_204[3:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (reset) begin
      wPos <= 6'h0;
    end else begin
      if (io_push) begin
        wPos <= _T_150;
      end
    end
    if (reset) begin
      rPos <= 3'h0;
    end else begin
      if (io_pop) begin
        rPos <= _T_153;
      end
    end
    if (io_push) begin
      if (6'h0 == wPos) begin
        mem_0 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h1 == wPos) begin
        mem_1 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h2 == wPos) begin
        mem_2 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h3 == wPos) begin
        mem_3 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h4 == wPos) begin
        mem_4 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h5 == wPos) begin
        mem_5 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h6 == wPos) begin
        mem_6 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h7 == wPos) begin
        mem_7 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h8 == wPos) begin
        mem_8 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h9 == wPos) begin
        mem_9 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'ha == wPos) begin
        mem_10 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'hb == wPos) begin
        mem_11 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'hc == wPos) begin
        mem_12 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'hd == wPos) begin
        mem_13 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'he == wPos) begin
        mem_14 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'hf == wPos) begin
        mem_15 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h10 == wPos) begin
        mem_16 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h11 == wPos) begin
        mem_17 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h12 == wPos) begin
        mem_18 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h13 == wPos) begin
        mem_19 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h14 == wPos) begin
        mem_20 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h15 == wPos) begin
        mem_21 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h16 == wPos) begin
        mem_22 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h17 == wPos) begin
        mem_23 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h18 == wPos) begin
        mem_24 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h19 == wPos) begin
        mem_25 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h1a == wPos) begin
        mem_26 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h1b == wPos) begin
        mem_27 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h1c == wPos) begin
        mem_28 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h1d == wPos) begin
        mem_29 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h1e == wPos) begin
        mem_30 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h1f == wPos) begin
        mem_31 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h20 == wPos) begin
        mem_32 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h21 == wPos) begin
        mem_33 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h22 == wPos) begin
        mem_34 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h23 == wPos) begin
        mem_35 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h24 == wPos) begin
        mem_36 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h25 == wPos) begin
        mem_37 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h26 == wPos) begin
        mem_38 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h27 == wPos) begin
        mem_39 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h28 == wPos) begin
        mem_40 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h29 == wPos) begin
        mem_41 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h2a == wPos) begin
        mem_42 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h2b == wPos) begin
        mem_43 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h2c == wPos) begin
        mem_44 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h2d == wPos) begin
        mem_45 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h2e == wPos) begin
        mem_46 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h2f == wPos) begin
        mem_47 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h30 == wPos) begin
        mem_48 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h31 == wPos) begin
        mem_49 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h32 == wPos) begin
        mem_50 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h33 == wPos) begin
        mem_51 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h34 == wPos) begin
        mem_52 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h35 == wPos) begin
        mem_53 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h36 == wPos) begin
        mem_54 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h37 == wPos) begin
        mem_55 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h38 == wPos) begin
        mem_56 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h39 == wPos) begin
        mem_57 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h3a == wPos) begin
        mem_58 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h3b == wPos) begin
        mem_59 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h3c == wPos) begin
        mem_60 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h3d == wPos) begin
        mem_61 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h3e == wPos) begin
        mem_62 <= _GEN_0;
      end
    end
    if (io_push) begin
      if (6'h3f == wPos) begin
        mem_63 <= _GEN_0;
      end
    end
  end
endmodule
module XNOR(
  input  [31:0] io_in1,
  input  [31:0] io_in2_0,
  input  [31:0] io_in2_1,
  input  [31:0] io_in2_2,
  input  [31:0] io_in2_3,
  output [31:0] io_out_0,
  output [31:0] io_out_1,
  output [31:0] io_out_2,
  output [31:0] io_out_3
);
  wire [31:0] _T_21;
  wire [31:0] _T_22;
  wire [31:0] _T_23;
  wire [31:0] _T_24;
  wire [31:0] _T_25;
  wire [31:0] _T_26;
  wire [31:0] _T_27;
  wire [31:0] _T_28;
  assign io_out_0 = _T_22;
  assign io_out_1 = _T_24;
  assign io_out_2 = _T_26;
  assign io_out_3 = _T_28;
  assign _T_21 = io_in1 ^ io_in2_0;
  assign _T_22 = ~ _T_21;
  assign _T_23 = io_in1 ^ io_in2_1;
  assign _T_24 = ~ _T_23;
  assign _T_25 = io_in1 ^ io_in2_2;
  assign _T_26 = ~ _T_25;
  assign _T_27 = io_in1 ^ io_in2_3;
  assign _T_28 = ~ _T_27;
endmodule
module MeanBuffer(
  input         clock,
  input         reset,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [15:0] io_cntInverse65536,
  input         io_reset,
  output [31:0] io_out
);
  reg [31:0] acc;
  reg [31:0] _GEN_3;
  wire  _T_17;
  wire [32:0] _T_19;
  wire [31:0] _T_20;
  wire [31:0] _T_21;
  wire [31:0] _T_22;
  wire [31:0] _T_23;
  wire  _T_25;
  wire [32:0] _T_27;
  wire [31:0] _T_28;
  wire [31:0] _T_29;
  wire [31:0] _T_30;
  wire [31:0] _T_31;
  wire  _T_33;
  wire [32:0] _T_35;
  wire [31:0] _T_36;
  wire [31:0] _T_37;
  wire [31:0] _T_38;
  wire [31:0] _T_39;
  wire  _T_41;
  wire [32:0] _T_43;
  wire [31:0] _T_44;
  wire [31:0] _T_45;
  wire [31:0] _T_46;
  wire [31:0] _T_47;
  wire [32:0] _T_48;
  wire [31:0] _T_49;
  wire [32:0] _T_50;
  wire [31:0] _T_51;
  wire [32:0] _T_52;
  wire [31:0] absSum;
  wire  _T_54;
  wire [32:0] _T_55;
  wire [31:0] _T_56;
  wire [31:0] _GEN_0;
  wire  _T_58;
  wire [31:0] _GEN_1;
  wire [31:0] _GEN_2;
  wire [47:0] _T_59;
  wire [31:0] _T_60;
  assign io_out = _T_60;
  assign _T_17 = $signed(io_in_0) > $signed(32'sh0);
  assign _T_19 = $signed(32'sh0) - $signed(io_in_0);
  assign _T_20 = _T_19[31:0];
  assign _T_21 = $signed(_T_20);
  assign _T_22 = _T_17 ? $signed(io_in_0) : $signed(_T_21);
  assign _T_23 = $unsigned(_T_22);
  assign _T_25 = $signed(io_in_1) > $signed(32'sh0);
  assign _T_27 = $signed(32'sh0) - $signed(io_in_1);
  assign _T_28 = _T_27[31:0];
  assign _T_29 = $signed(_T_28);
  assign _T_30 = _T_25 ? $signed(io_in_1) : $signed(_T_29);
  assign _T_31 = $unsigned(_T_30);
  assign _T_33 = $signed(io_in_2) > $signed(32'sh0);
  assign _T_35 = $signed(32'sh0) - $signed(io_in_2);
  assign _T_36 = _T_35[31:0];
  assign _T_37 = $signed(_T_36);
  assign _T_38 = _T_33 ? $signed(io_in_2) : $signed(_T_37);
  assign _T_39 = $unsigned(_T_38);
  assign _T_41 = $signed(io_in_3) > $signed(32'sh0);
  assign _T_43 = $signed(32'sh0) - $signed(io_in_3);
  assign _T_44 = _T_43[31:0];
  assign _T_45 = $signed(_T_44);
  assign _T_46 = _T_41 ? $signed(io_in_3) : $signed(_T_45);
  assign _T_47 = $unsigned(_T_46);
  assign _T_48 = _T_23 + _T_31;
  assign _T_49 = _T_48[31:0];
  assign _T_50 = _T_39 + _T_47;
  assign _T_51 = _T_50[31:0];
  assign _T_52 = _T_49 + _T_51;
  assign absSum = _T_52[31:0];
  assign _T_54 = io_reset == 1'h0;
  assign _T_55 = acc + absSum;
  assign _T_56 = _T_55[31:0];
  assign _GEN_0 = _T_54 ? _T_56 : acc;
  assign _T_58 = _T_54 == 1'h0;
  assign _GEN_1 = _T_58 ? absSum : _GEN_0;
  assign _GEN_2 = {{16'd0}, io_cntInverse65536};
  assign _T_59 = acc * _GEN_2;
  assign _T_60 = _T_59[47:16];
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_3 = {1{$random}};
  acc = _GEN_3[31:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (reset) begin
      acc <= 32'h0;
    end else begin
      if (_T_58) begin
        acc <= absSum;
      end else begin
        if (_T_54) begin
          acc <= _T_56;
        end
      end
    end
  end
endmodule
module DelayedOutput(
  input         clock,
  input         reset,
  input  [31:0] io_input,
  input         io_update,
  output [31:0] io_output
);
  reg [31:0] reg$;
  reg [31:0] _GEN_1;
  wire [31:0] _GEN_0;
  assign io_output = reg$;
  assign _GEN_0 = io_update ? io_input : reg$;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1 = {1{$random}};
  reg$ = _GEN_1[31:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (reset) begin
      reg$ <= 32'h1;
    end else begin
      if (io_update) begin
        reg$ <= io_input;
      end
    end
  end
endmodule
module MaxBuffer(
  input         clock,
  input         io_reset,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [3:0]  io_offset,
  output [3:0]  io_out
);
  reg [3:0] idxReg;
  reg [31:0] _GEN_6;
  reg [31:0] dataReg;
  reg [31:0] _GEN_7;
  wire [4:0] _T_18;
  wire [3:0] _T_19;
  wire [4:0] _T_21;
  wire [3:0] _T_22;
  wire [4:0] _T_24;
  wire [3:0] _T_25;
  wire [4:0] _T_27;
  wire [3:0] _T_28;
  wire  _T_29;
  wire [3:0] _T_30;
  wire [31:0] _T_31;
  wire  _T_32;
  wire [3:0] _T_33;
  wire [31:0] _T_34;
  wire  _T_35;
  wire [3:0] _T_36;
  wire [31:0] _T_37;
  wire  cmp2;
  wire  _T_39;
  wire [31:0] _T_40;
  wire [3:0] _T_41;
  wire [31:0] _GEN_0;
  wire [3:0] _GEN_1;
  wire  _T_43;
  wire [31:0] _GEN_2;
  wire [3:0] _GEN_3;
  wire [31:0] _GEN_4;
  wire [3:0] _GEN_5;
  assign io_out = idxReg;
  assign _T_18 = 4'h0 + io_offset;
  assign _T_19 = _T_18[3:0];
  assign _T_21 = 4'h1 + io_offset;
  assign _T_22 = _T_21[3:0];
  assign _T_24 = 4'h2 + io_offset;
  assign _T_25 = _T_24[3:0];
  assign _T_27 = 4'h3 + io_offset;
  assign _T_28 = _T_27[3:0];
  assign _T_29 = $signed(io_in_0) > $signed(io_in_1);
  assign _T_30 = _T_29 ? _T_19 : _T_22;
  assign _T_31 = _T_29 ? $signed(io_in_0) : $signed(io_in_1);
  assign _T_32 = $signed(io_in_2) > $signed(io_in_3);
  assign _T_33 = _T_32 ? _T_25 : _T_28;
  assign _T_34 = _T_32 ? $signed(io_in_2) : $signed(io_in_3);
  assign _T_35 = $signed(_T_31) > $signed(_T_34);
  assign _T_36 = _T_35 ? _T_30 : _T_33;
  assign _T_37 = _T_35 ? $signed(_T_31) : $signed(_T_34);
  assign cmp2 = $signed(dataReg) > $signed(_T_37);
  assign _T_39 = io_reset == 1'h0;
  assign _T_40 = cmp2 ? $signed(dataReg) : $signed(_T_37);
  assign _T_41 = cmp2 ? idxReg : _T_36;
  assign _GEN_0 = _T_39 ? $signed(_T_40) : $signed(dataReg);
  assign _GEN_1 = _T_39 ? _T_41 : idxReg;
  assign _T_43 = _T_39 == 1'h0;
  assign _GEN_2 = _T_43 ? $signed(_T_37) : $signed(_GEN_0);
  assign _GEN_3 = _T_43 ? _T_36 : _GEN_1;
  assign _GEN_4 = io_en ? $signed(_GEN_2) : $signed(dataReg);
  assign _GEN_5 = io_en ? _GEN_3 : idxReg;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_6 = {1{$random}};
  idxReg = _GEN_6[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_7 = {1{$random}};
  dataReg = _GEN_7[31:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (io_en) begin
      if (_T_43) begin
        if (_T_35) begin
          if (_T_29) begin
            idxReg <= _T_19;
          end else begin
            idxReg <= _T_22;
          end
        end else begin
          if (_T_32) begin
            idxReg <= _T_25;
          end else begin
            idxReg <= _T_28;
          end
        end
      end else begin
        if (_T_39) begin
          if (!(cmp2)) begin
            if (_T_35) begin
              if (_T_29) begin
                idxReg <= _T_19;
              end else begin
                idxReg <= _T_22;
              end
            end else begin
              if (_T_32) begin
                idxReg <= _T_25;
              end else begin
                idxReg <= _T_28;
              end
            end
          end
        end
      end
    end
    if (io_en) begin
      if (_T_43) begin
        if (_T_35) begin
          if (_T_29) begin
            dataReg <= io_in_0;
          end else begin
            dataReg <= io_in_1;
          end
        end else begin
          if (_T_32) begin
            dataReg <= io_in_2;
          end else begin
            dataReg <= io_in_3;
          end
        end
      end else begin
        if (_T_39) begin
          if (!(cmp2)) begin
            if (_T_35) begin
              if (_T_29) begin
                dataReg <= io_in_0;
              end else begin
                dataReg <= io_in_1;
              end
            end else begin
              if (_T_32) begin
                dataReg <= io_in_2;
              end else begin
                dataReg <= io_in_3;
              end
            end
          end
        end
      end
    end
  end
endmodule
module Accumulator(
  input         clock,
  input  [31:0] io_in,
  output [31:0] io_out,
  input  [4:0]  io_sel,
  input         io_en,
  input         io_reset
);
  reg [31:0] accumulator_0;
  reg [31:0] _GEN_131;
  reg [31:0] accumulator_1;
  reg [31:0] _GEN_132;
  reg [31:0] accumulator_2;
  reg [31:0] _GEN_133;
  reg [31:0] accumulator_3;
  reg [31:0] _GEN_134;
  reg [31:0] accumulator_4;
  reg [31:0] _GEN_135;
  reg [31:0] accumulator_5;
  reg [31:0] _GEN_136;
  reg [31:0] accumulator_6;
  reg [31:0] _GEN_137;
  reg [31:0] accumulator_7;
  reg [31:0] _GEN_138;
  reg [31:0] accumulator_8;
  reg [31:0] _GEN_139;
  reg [31:0] accumulator_9;
  reg [31:0] _GEN_140;
  reg [31:0] accumulator_10;
  reg [31:0] _GEN_141;
  reg [31:0] accumulator_11;
  reg [31:0] _GEN_142;
  reg [31:0] accumulator_12;
  reg [31:0] _GEN_143;
  reg [31:0] accumulator_13;
  reg [31:0] _GEN_144;
  reg [31:0] accumulator_14;
  reg [31:0] _GEN_145;
  reg [31:0] accumulator_15;
  reg [31:0] _GEN_146;
  reg [31:0] accumulator_16;
  reg [31:0] _GEN_147;
  reg [31:0] accumulator_17;
  reg [31:0] _GEN_148;
  reg [31:0] accumulator_18;
  reg [31:0] _GEN_149;
  reg [31:0] accumulator_19;
  reg [31:0] _GEN_150;
  reg [31:0] accumulator_20;
  reg [31:0] _GEN_151;
  reg [31:0] accumulator_21;
  reg [31:0] _GEN_152;
  reg [31:0] accumulator_22;
  reg [31:0] _GEN_153;
  reg [31:0] accumulator_23;
  reg [31:0] _GEN_154;
  reg [31:0] accumulator_24;
  reg [31:0] _GEN_155;
  reg [31:0] accumulator_25;
  reg [31:0] _GEN_156;
  reg [31:0] accumulator_26;
  reg [31:0] _GEN_157;
  reg [31:0] accumulator_27;
  reg [31:0] _GEN_158;
  reg [31:0] accumulator_28;
  reg [31:0] _GEN_159;
  reg [31:0] accumulator_29;
  reg [31:0] _GEN_160;
  reg [31:0] accumulator_30;
  reg [31:0] _GEN_161;
  reg [31:0] accumulator_31;
  reg [31:0] _GEN_162;
  wire  _T_46;
  wire  _T_47;
  wire [31:0] _GEN_0;
  wire [31:0] _GEN_3;
  wire [31:0] _GEN_4;
  wire [31:0] _GEN_5;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_7;
  wire [31:0] _GEN_8;
  wire [31:0] _GEN_9;
  wire [31:0] _GEN_10;
  wire [31:0] _GEN_11;
  wire [31:0] _GEN_12;
  wire [31:0] _GEN_13;
  wire [31:0] _GEN_14;
  wire [31:0] _GEN_15;
  wire [31:0] _GEN_16;
  wire [31:0] _GEN_17;
  wire [31:0] _GEN_18;
  wire [31:0] _GEN_19;
  wire [31:0] _GEN_20;
  wire [31:0] _GEN_21;
  wire [31:0] _GEN_22;
  wire [31:0] _GEN_23;
  wire [31:0] _GEN_24;
  wire [31:0] _GEN_25;
  wire [31:0] _GEN_26;
  wire [31:0] _GEN_27;
  wire [31:0] _GEN_28;
  wire [31:0] _GEN_29;
  wire [31:0] _GEN_30;
  wire [31:0] _GEN_31;
  wire [31:0] _GEN_32;
  wire [31:0] _GEN_33;
  wire [32:0] _T_48;
  wire [31:0] _T_49;
  wire [31:0] _T_50;
  wire [31:0] _GEN_1;
  wire [31:0] _GEN_34;
  wire [31:0] _GEN_35;
  wire [31:0] _GEN_36;
  wire [31:0] _GEN_37;
  wire [31:0] _GEN_38;
  wire [31:0] _GEN_39;
  wire [31:0] _GEN_40;
  wire [31:0] _GEN_41;
  wire [31:0] _GEN_42;
  wire [31:0] _GEN_43;
  wire [31:0] _GEN_44;
  wire [31:0] _GEN_45;
  wire [31:0] _GEN_46;
  wire [31:0] _GEN_47;
  wire [31:0] _GEN_48;
  wire [31:0] _GEN_49;
  wire [31:0] _GEN_50;
  wire [31:0] _GEN_51;
  wire [31:0] _GEN_52;
  wire [31:0] _GEN_53;
  wire [31:0] _GEN_54;
  wire [31:0] _GEN_55;
  wire [31:0] _GEN_56;
  wire [31:0] _GEN_57;
  wire [31:0] _GEN_58;
  wire [31:0] _GEN_59;
  wire [31:0] _GEN_60;
  wire [31:0] _GEN_61;
  wire [31:0] _GEN_62;
  wire [31:0] _GEN_63;
  wire [31:0] _GEN_64;
  wire [31:0] _GEN_65;
  wire [31:0] _GEN_66;
  wire [31:0] _GEN_67;
  wire [31:0] _GEN_68;
  wire [31:0] _GEN_69;
  wire [31:0] _GEN_70;
  wire [31:0] _GEN_71;
  wire [31:0] _GEN_72;
  wire [31:0] _GEN_73;
  wire [31:0] _GEN_74;
  wire [31:0] _GEN_75;
  wire [31:0] _GEN_76;
  wire [31:0] _GEN_77;
  wire [31:0] _GEN_78;
  wire [31:0] _GEN_79;
  wire [31:0] _GEN_80;
  wire [31:0] _GEN_81;
  wire [31:0] _GEN_82;
  wire [31:0] _GEN_83;
  wire [31:0] _GEN_84;
  wire [31:0] _GEN_85;
  wire [31:0] _GEN_86;
  wire [31:0] _GEN_87;
  wire [31:0] _GEN_88;
  wire [31:0] _GEN_89;
  wire [31:0] _GEN_90;
  wire [31:0] _GEN_91;
  wire [31:0] _GEN_92;
  wire [31:0] _GEN_93;
  wire [31:0] _GEN_94;
  wire [31:0] _GEN_95;
  wire [31:0] _GEN_96;
  wire [31:0] _GEN_97;
  wire [31:0] _GEN_2;
  wire  _T_51;
  wire  _T_53;
  wire [31:0] _T_55;
  wire  _T_57;
  wire [31:0] _T_59;
  wire  _T_61;
  wire [31:0] _T_63;
  wire  _T_65;
  wire [31:0] _T_67;
  wire  _T_69;
  wire [31:0] _T_71;
  wire  _T_73;
  wire [31:0] _T_75;
  wire  _T_77;
  wire [31:0] _T_79;
  wire  _T_81;
  wire [31:0] _T_83;
  wire  _T_85;
  wire [31:0] _T_87;
  wire  _T_89;
  wire [31:0] _T_91;
  wire  _T_93;
  wire [31:0] _T_95;
  wire  _T_97;
  wire [31:0] _T_99;
  wire  _T_101;
  wire [31:0] _T_103;
  wire  _T_105;
  wire [31:0] _T_107;
  wire  _T_109;
  wire [31:0] _T_111;
  wire  _T_113;
  wire [31:0] _T_115;
  wire  _T_117;
  wire [31:0] _T_119;
  wire  _T_121;
  wire [31:0] _T_123;
  wire  _T_125;
  wire [31:0] _T_127;
  wire  _T_129;
  wire [31:0] _T_131;
  wire  _T_133;
  wire [31:0] _T_135;
  wire  _T_137;
  wire [31:0] _T_139;
  wire  _T_141;
  wire [31:0] _T_143;
  wire  _T_145;
  wire [31:0] _T_147;
  wire  _T_149;
  wire [31:0] _T_151;
  wire  _T_153;
  wire [31:0] _T_155;
  wire  _T_157;
  wire [31:0] _T_159;
  wire  _T_161;
  wire [31:0] _T_163;
  wire  _T_165;
  wire [31:0] _T_167;
  wire  _T_169;
  wire [31:0] _T_171;
  wire  _T_173;
  wire [31:0] _T_175;
  wire  _T_177;
  wire [31:0] _T_179;
  wire [31:0] _GEN_98;
  wire [31:0] _GEN_99;
  wire [31:0] _GEN_100;
  wire [31:0] _GEN_101;
  wire [31:0] _GEN_102;
  wire [31:0] _GEN_103;
  wire [31:0] _GEN_104;
  wire [31:0] _GEN_105;
  wire [31:0] _GEN_106;
  wire [31:0] _GEN_107;
  wire [31:0] _GEN_108;
  wire [31:0] _GEN_109;
  wire [31:0] _GEN_110;
  wire [31:0] _GEN_111;
  wire [31:0] _GEN_112;
  wire [31:0] _GEN_113;
  wire [31:0] _GEN_114;
  wire [31:0] _GEN_115;
  wire [31:0] _GEN_116;
  wire [31:0] _GEN_117;
  wire [31:0] _GEN_118;
  wire [31:0] _GEN_119;
  wire [31:0] _GEN_120;
  wire [31:0] _GEN_121;
  wire [31:0] _GEN_122;
  wire [31:0] _GEN_123;
  wire [31:0] _GEN_124;
  wire [31:0] _GEN_125;
  wire [31:0] _GEN_126;
  wire [31:0] _GEN_127;
  wire [31:0] _GEN_128;
  wire [31:0] _GEN_129;
  wire [31:0] _GEN_130;
  assign io_out = _GEN_130;
  assign _T_46 = io_reset == 1'h0;
  assign _T_47 = io_en & _T_46;
  assign _GEN_0 = _GEN_33;
  assign _GEN_3 = 5'h1 == io_sel ? $signed(accumulator_1) : $signed(accumulator_0);
  assign _GEN_4 = 5'h2 == io_sel ? $signed(accumulator_2) : $signed(_GEN_3);
  assign _GEN_5 = 5'h3 == io_sel ? $signed(accumulator_3) : $signed(_GEN_4);
  assign _GEN_6 = 5'h4 == io_sel ? $signed(accumulator_4) : $signed(_GEN_5);
  assign _GEN_7 = 5'h5 == io_sel ? $signed(accumulator_5) : $signed(_GEN_6);
  assign _GEN_8 = 5'h6 == io_sel ? $signed(accumulator_6) : $signed(_GEN_7);
  assign _GEN_9 = 5'h7 == io_sel ? $signed(accumulator_7) : $signed(_GEN_8);
  assign _GEN_10 = 5'h8 == io_sel ? $signed(accumulator_8) : $signed(_GEN_9);
  assign _GEN_11 = 5'h9 == io_sel ? $signed(accumulator_9) : $signed(_GEN_10);
  assign _GEN_12 = 5'ha == io_sel ? $signed(accumulator_10) : $signed(_GEN_11);
  assign _GEN_13 = 5'hb == io_sel ? $signed(accumulator_11) : $signed(_GEN_12);
  assign _GEN_14 = 5'hc == io_sel ? $signed(accumulator_12) : $signed(_GEN_13);
  assign _GEN_15 = 5'hd == io_sel ? $signed(accumulator_13) : $signed(_GEN_14);
  assign _GEN_16 = 5'he == io_sel ? $signed(accumulator_14) : $signed(_GEN_15);
  assign _GEN_17 = 5'hf == io_sel ? $signed(accumulator_15) : $signed(_GEN_16);
  assign _GEN_18 = 5'h10 == io_sel ? $signed(accumulator_16) : $signed(_GEN_17);
  assign _GEN_19 = 5'h11 == io_sel ? $signed(accumulator_17) : $signed(_GEN_18);
  assign _GEN_20 = 5'h12 == io_sel ? $signed(accumulator_18) : $signed(_GEN_19);
  assign _GEN_21 = 5'h13 == io_sel ? $signed(accumulator_19) : $signed(_GEN_20);
  assign _GEN_22 = 5'h14 == io_sel ? $signed(accumulator_20) : $signed(_GEN_21);
  assign _GEN_23 = 5'h15 == io_sel ? $signed(accumulator_21) : $signed(_GEN_22);
  assign _GEN_24 = 5'h16 == io_sel ? $signed(accumulator_22) : $signed(_GEN_23);
  assign _GEN_25 = 5'h17 == io_sel ? $signed(accumulator_23) : $signed(_GEN_24);
  assign _GEN_26 = 5'h18 == io_sel ? $signed(accumulator_24) : $signed(_GEN_25);
  assign _GEN_27 = 5'h19 == io_sel ? $signed(accumulator_25) : $signed(_GEN_26);
  assign _GEN_28 = 5'h1a == io_sel ? $signed(accumulator_26) : $signed(_GEN_27);
  assign _GEN_29 = 5'h1b == io_sel ? $signed(accumulator_27) : $signed(_GEN_28);
  assign _GEN_30 = 5'h1c == io_sel ? $signed(accumulator_28) : $signed(_GEN_29);
  assign _GEN_31 = 5'h1d == io_sel ? $signed(accumulator_29) : $signed(_GEN_30);
  assign _GEN_32 = 5'h1e == io_sel ? $signed(accumulator_30) : $signed(_GEN_31);
  assign _GEN_33 = 5'h1f == io_sel ? $signed(accumulator_31) : $signed(_GEN_32);
  assign _T_48 = $signed(_GEN_0) + $signed(io_in);
  assign _T_49 = _T_48[31:0];
  assign _T_50 = $signed(_T_49);
  assign _GEN_1 = _T_50;
  assign _GEN_34 = 5'h0 == io_sel ? $signed(_GEN_1) : $signed(accumulator_0);
  assign _GEN_35 = 5'h1 == io_sel ? $signed(_GEN_1) : $signed(accumulator_1);
  assign _GEN_36 = 5'h2 == io_sel ? $signed(_GEN_1) : $signed(accumulator_2);
  assign _GEN_37 = 5'h3 == io_sel ? $signed(_GEN_1) : $signed(accumulator_3);
  assign _GEN_38 = 5'h4 == io_sel ? $signed(_GEN_1) : $signed(accumulator_4);
  assign _GEN_39 = 5'h5 == io_sel ? $signed(_GEN_1) : $signed(accumulator_5);
  assign _GEN_40 = 5'h6 == io_sel ? $signed(_GEN_1) : $signed(accumulator_6);
  assign _GEN_41 = 5'h7 == io_sel ? $signed(_GEN_1) : $signed(accumulator_7);
  assign _GEN_42 = 5'h8 == io_sel ? $signed(_GEN_1) : $signed(accumulator_8);
  assign _GEN_43 = 5'h9 == io_sel ? $signed(_GEN_1) : $signed(accumulator_9);
  assign _GEN_44 = 5'ha == io_sel ? $signed(_GEN_1) : $signed(accumulator_10);
  assign _GEN_45 = 5'hb == io_sel ? $signed(_GEN_1) : $signed(accumulator_11);
  assign _GEN_46 = 5'hc == io_sel ? $signed(_GEN_1) : $signed(accumulator_12);
  assign _GEN_47 = 5'hd == io_sel ? $signed(_GEN_1) : $signed(accumulator_13);
  assign _GEN_48 = 5'he == io_sel ? $signed(_GEN_1) : $signed(accumulator_14);
  assign _GEN_49 = 5'hf == io_sel ? $signed(_GEN_1) : $signed(accumulator_15);
  assign _GEN_50 = 5'h10 == io_sel ? $signed(_GEN_1) : $signed(accumulator_16);
  assign _GEN_51 = 5'h11 == io_sel ? $signed(_GEN_1) : $signed(accumulator_17);
  assign _GEN_52 = 5'h12 == io_sel ? $signed(_GEN_1) : $signed(accumulator_18);
  assign _GEN_53 = 5'h13 == io_sel ? $signed(_GEN_1) : $signed(accumulator_19);
  assign _GEN_54 = 5'h14 == io_sel ? $signed(_GEN_1) : $signed(accumulator_20);
  assign _GEN_55 = 5'h15 == io_sel ? $signed(_GEN_1) : $signed(accumulator_21);
  assign _GEN_56 = 5'h16 == io_sel ? $signed(_GEN_1) : $signed(accumulator_22);
  assign _GEN_57 = 5'h17 == io_sel ? $signed(_GEN_1) : $signed(accumulator_23);
  assign _GEN_58 = 5'h18 == io_sel ? $signed(_GEN_1) : $signed(accumulator_24);
  assign _GEN_59 = 5'h19 == io_sel ? $signed(_GEN_1) : $signed(accumulator_25);
  assign _GEN_60 = 5'h1a == io_sel ? $signed(_GEN_1) : $signed(accumulator_26);
  assign _GEN_61 = 5'h1b == io_sel ? $signed(_GEN_1) : $signed(accumulator_27);
  assign _GEN_62 = 5'h1c == io_sel ? $signed(_GEN_1) : $signed(accumulator_28);
  assign _GEN_63 = 5'h1d == io_sel ? $signed(_GEN_1) : $signed(accumulator_29);
  assign _GEN_64 = 5'h1e == io_sel ? $signed(_GEN_1) : $signed(accumulator_30);
  assign _GEN_65 = 5'h1f == io_sel ? $signed(_GEN_1) : $signed(accumulator_31);
  assign _GEN_66 = _T_47 ? $signed(_GEN_34) : $signed(accumulator_0);
  assign _GEN_67 = _T_47 ? $signed(_GEN_35) : $signed(accumulator_1);
  assign _GEN_68 = _T_47 ? $signed(_GEN_36) : $signed(accumulator_2);
  assign _GEN_69 = _T_47 ? $signed(_GEN_37) : $signed(accumulator_3);
  assign _GEN_70 = _T_47 ? $signed(_GEN_38) : $signed(accumulator_4);
  assign _GEN_71 = _T_47 ? $signed(_GEN_39) : $signed(accumulator_5);
  assign _GEN_72 = _T_47 ? $signed(_GEN_40) : $signed(accumulator_6);
  assign _GEN_73 = _T_47 ? $signed(_GEN_41) : $signed(accumulator_7);
  assign _GEN_74 = _T_47 ? $signed(_GEN_42) : $signed(accumulator_8);
  assign _GEN_75 = _T_47 ? $signed(_GEN_43) : $signed(accumulator_9);
  assign _GEN_76 = _T_47 ? $signed(_GEN_44) : $signed(accumulator_10);
  assign _GEN_77 = _T_47 ? $signed(_GEN_45) : $signed(accumulator_11);
  assign _GEN_78 = _T_47 ? $signed(_GEN_46) : $signed(accumulator_12);
  assign _GEN_79 = _T_47 ? $signed(_GEN_47) : $signed(accumulator_13);
  assign _GEN_80 = _T_47 ? $signed(_GEN_48) : $signed(accumulator_14);
  assign _GEN_81 = _T_47 ? $signed(_GEN_49) : $signed(accumulator_15);
  assign _GEN_82 = _T_47 ? $signed(_GEN_50) : $signed(accumulator_16);
  assign _GEN_83 = _T_47 ? $signed(_GEN_51) : $signed(accumulator_17);
  assign _GEN_84 = _T_47 ? $signed(_GEN_52) : $signed(accumulator_18);
  assign _GEN_85 = _T_47 ? $signed(_GEN_53) : $signed(accumulator_19);
  assign _GEN_86 = _T_47 ? $signed(_GEN_54) : $signed(accumulator_20);
  assign _GEN_87 = _T_47 ? $signed(_GEN_55) : $signed(accumulator_21);
  assign _GEN_88 = _T_47 ? $signed(_GEN_56) : $signed(accumulator_22);
  assign _GEN_89 = _T_47 ? $signed(_GEN_57) : $signed(accumulator_23);
  assign _GEN_90 = _T_47 ? $signed(_GEN_58) : $signed(accumulator_24);
  assign _GEN_91 = _T_47 ? $signed(_GEN_59) : $signed(accumulator_25);
  assign _GEN_92 = _T_47 ? $signed(_GEN_60) : $signed(accumulator_26);
  assign _GEN_93 = _T_47 ? $signed(_GEN_61) : $signed(accumulator_27);
  assign _GEN_94 = _T_47 ? $signed(_GEN_62) : $signed(accumulator_28);
  assign _GEN_95 = _T_47 ? $signed(_GEN_63) : $signed(accumulator_29);
  assign _GEN_96 = _T_47 ? $signed(_GEN_64) : $signed(accumulator_30);
  assign _GEN_97 = _T_47 ? $signed(_GEN_65) : $signed(accumulator_31);
  assign _GEN_2 = _GEN_33;
  assign _T_51 = io_en & io_reset;
  assign _T_53 = 5'h0 == io_sel;
  assign _T_55 = _T_53 ? $signed(io_in) : $signed(32'sh0);
  assign _T_57 = 5'h1 == io_sel;
  assign _T_59 = _T_57 ? $signed(io_in) : $signed(32'sh0);
  assign _T_61 = 5'h2 == io_sel;
  assign _T_63 = _T_61 ? $signed(io_in) : $signed(32'sh0);
  assign _T_65 = 5'h3 == io_sel;
  assign _T_67 = _T_65 ? $signed(io_in) : $signed(32'sh0);
  assign _T_69 = 5'h4 == io_sel;
  assign _T_71 = _T_69 ? $signed(io_in) : $signed(32'sh0);
  assign _T_73 = 5'h5 == io_sel;
  assign _T_75 = _T_73 ? $signed(io_in) : $signed(32'sh0);
  assign _T_77 = 5'h6 == io_sel;
  assign _T_79 = _T_77 ? $signed(io_in) : $signed(32'sh0);
  assign _T_81 = 5'h7 == io_sel;
  assign _T_83 = _T_81 ? $signed(io_in) : $signed(32'sh0);
  assign _T_85 = 5'h8 == io_sel;
  assign _T_87 = _T_85 ? $signed(io_in) : $signed(32'sh0);
  assign _T_89 = 5'h9 == io_sel;
  assign _T_91 = _T_89 ? $signed(io_in) : $signed(32'sh0);
  assign _T_93 = 5'ha == io_sel;
  assign _T_95 = _T_93 ? $signed(io_in) : $signed(32'sh0);
  assign _T_97 = 5'hb == io_sel;
  assign _T_99 = _T_97 ? $signed(io_in) : $signed(32'sh0);
  assign _T_101 = 5'hc == io_sel;
  assign _T_103 = _T_101 ? $signed(io_in) : $signed(32'sh0);
  assign _T_105 = 5'hd == io_sel;
  assign _T_107 = _T_105 ? $signed(io_in) : $signed(32'sh0);
  assign _T_109 = 5'he == io_sel;
  assign _T_111 = _T_109 ? $signed(io_in) : $signed(32'sh0);
  assign _T_113 = 5'hf == io_sel;
  assign _T_115 = _T_113 ? $signed(io_in) : $signed(32'sh0);
  assign _T_117 = 5'h10 == io_sel;
  assign _T_119 = _T_117 ? $signed(io_in) : $signed(32'sh0);
  assign _T_121 = 5'h11 == io_sel;
  assign _T_123 = _T_121 ? $signed(io_in) : $signed(32'sh0);
  assign _T_125 = 5'h12 == io_sel;
  assign _T_127 = _T_125 ? $signed(io_in) : $signed(32'sh0);
  assign _T_129 = 5'h13 == io_sel;
  assign _T_131 = _T_129 ? $signed(io_in) : $signed(32'sh0);
  assign _T_133 = 5'h14 == io_sel;
  assign _T_135 = _T_133 ? $signed(io_in) : $signed(32'sh0);
  assign _T_137 = 5'h15 == io_sel;
  assign _T_139 = _T_137 ? $signed(io_in) : $signed(32'sh0);
  assign _T_141 = 5'h16 == io_sel;
  assign _T_143 = _T_141 ? $signed(io_in) : $signed(32'sh0);
  assign _T_145 = 5'h17 == io_sel;
  assign _T_147 = _T_145 ? $signed(io_in) : $signed(32'sh0);
  assign _T_149 = 5'h18 == io_sel;
  assign _T_151 = _T_149 ? $signed(io_in) : $signed(32'sh0);
  assign _T_153 = 5'h19 == io_sel;
  assign _T_155 = _T_153 ? $signed(io_in) : $signed(32'sh0);
  assign _T_157 = 5'h1a == io_sel;
  assign _T_159 = _T_157 ? $signed(io_in) : $signed(32'sh0);
  assign _T_161 = 5'h1b == io_sel;
  assign _T_163 = _T_161 ? $signed(io_in) : $signed(32'sh0);
  assign _T_165 = 5'h1c == io_sel;
  assign _T_167 = _T_165 ? $signed(io_in) : $signed(32'sh0);
  assign _T_169 = 5'h1d == io_sel;
  assign _T_171 = _T_169 ? $signed(io_in) : $signed(32'sh0);
  assign _T_173 = 5'h1e == io_sel;
  assign _T_175 = _T_173 ? $signed(io_in) : $signed(32'sh0);
  assign _T_177 = 5'h1f == io_sel;
  assign _T_179 = _T_177 ? $signed(io_in) : $signed(32'sh0);
  assign _GEN_98 = _T_51 ? $signed(_T_55) : $signed(_GEN_66);
  assign _GEN_99 = _T_51 ? $signed(_T_59) : $signed(_GEN_67);
  assign _GEN_100 = _T_51 ? $signed(_T_63) : $signed(_GEN_68);
  assign _GEN_101 = _T_51 ? $signed(_T_67) : $signed(_GEN_69);
  assign _GEN_102 = _T_51 ? $signed(_T_71) : $signed(_GEN_70);
  assign _GEN_103 = _T_51 ? $signed(_T_75) : $signed(_GEN_71);
  assign _GEN_104 = _T_51 ? $signed(_T_79) : $signed(_GEN_72);
  assign _GEN_105 = _T_51 ? $signed(_T_83) : $signed(_GEN_73);
  assign _GEN_106 = _T_51 ? $signed(_T_87) : $signed(_GEN_74);
  assign _GEN_107 = _T_51 ? $signed(_T_91) : $signed(_GEN_75);
  assign _GEN_108 = _T_51 ? $signed(_T_95) : $signed(_GEN_76);
  assign _GEN_109 = _T_51 ? $signed(_T_99) : $signed(_GEN_77);
  assign _GEN_110 = _T_51 ? $signed(_T_103) : $signed(_GEN_78);
  assign _GEN_111 = _T_51 ? $signed(_T_107) : $signed(_GEN_79);
  assign _GEN_112 = _T_51 ? $signed(_T_111) : $signed(_GEN_80);
  assign _GEN_113 = _T_51 ? $signed(_T_115) : $signed(_GEN_81);
  assign _GEN_114 = _T_51 ? $signed(_T_119) : $signed(_GEN_82);
  assign _GEN_115 = _T_51 ? $signed(_T_123) : $signed(_GEN_83);
  assign _GEN_116 = _T_51 ? $signed(_T_127) : $signed(_GEN_84);
  assign _GEN_117 = _T_51 ? $signed(_T_131) : $signed(_GEN_85);
  assign _GEN_118 = _T_51 ? $signed(_T_135) : $signed(_GEN_86);
  assign _GEN_119 = _T_51 ? $signed(_T_139) : $signed(_GEN_87);
  assign _GEN_120 = _T_51 ? $signed(_T_143) : $signed(_GEN_88);
  assign _GEN_121 = _T_51 ? $signed(_T_147) : $signed(_GEN_89);
  assign _GEN_122 = _T_51 ? $signed(_T_151) : $signed(_GEN_90);
  assign _GEN_123 = _T_51 ? $signed(_T_155) : $signed(_GEN_91);
  assign _GEN_124 = _T_51 ? $signed(_T_159) : $signed(_GEN_92);
  assign _GEN_125 = _T_51 ? $signed(_T_163) : $signed(_GEN_93);
  assign _GEN_126 = _T_51 ? $signed(_T_167) : $signed(_GEN_94);
  assign _GEN_127 = _T_51 ? $signed(_T_171) : $signed(_GEN_95);
  assign _GEN_128 = _T_51 ? $signed(_T_175) : $signed(_GEN_96);
  assign _GEN_129 = _T_51 ? $signed(_T_179) : $signed(_GEN_97);
  assign _GEN_130 = _T_51 ? $signed(io_in) : $signed(_GEN_2);
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_131 = {1{$random}};
  accumulator_0 = _GEN_131[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_132 = {1{$random}};
  accumulator_1 = _GEN_132[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_133 = {1{$random}};
  accumulator_2 = _GEN_133[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_134 = {1{$random}};
  accumulator_3 = _GEN_134[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_135 = {1{$random}};
  accumulator_4 = _GEN_135[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_136 = {1{$random}};
  accumulator_5 = _GEN_136[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_137 = {1{$random}};
  accumulator_6 = _GEN_137[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_138 = {1{$random}};
  accumulator_7 = _GEN_138[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_139 = {1{$random}};
  accumulator_8 = _GEN_139[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_140 = {1{$random}};
  accumulator_9 = _GEN_140[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_141 = {1{$random}};
  accumulator_10 = _GEN_141[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_142 = {1{$random}};
  accumulator_11 = _GEN_142[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_143 = {1{$random}};
  accumulator_12 = _GEN_143[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_144 = {1{$random}};
  accumulator_13 = _GEN_144[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_145 = {1{$random}};
  accumulator_14 = _GEN_145[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_146 = {1{$random}};
  accumulator_15 = _GEN_146[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_147 = {1{$random}};
  accumulator_16 = _GEN_147[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_148 = {1{$random}};
  accumulator_17 = _GEN_148[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_149 = {1{$random}};
  accumulator_18 = _GEN_149[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_150 = {1{$random}};
  accumulator_19 = _GEN_150[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_151 = {1{$random}};
  accumulator_20 = _GEN_151[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_152 = {1{$random}};
  accumulator_21 = _GEN_152[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_153 = {1{$random}};
  accumulator_22 = _GEN_153[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_154 = {1{$random}};
  accumulator_23 = _GEN_154[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_155 = {1{$random}};
  accumulator_24 = _GEN_155[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_156 = {1{$random}};
  accumulator_25 = _GEN_156[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_157 = {1{$random}};
  accumulator_26 = _GEN_157[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_158 = {1{$random}};
  accumulator_27 = _GEN_158[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_159 = {1{$random}};
  accumulator_28 = _GEN_159[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_160 = {1{$random}};
  accumulator_29 = _GEN_160[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_161 = {1{$random}};
  accumulator_30 = _GEN_161[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_162 = {1{$random}};
  accumulator_31 = _GEN_162[31:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (_T_51) begin
      if (_T_53) begin
        accumulator_0 <= io_in;
      end else begin
        accumulator_0 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h0 == io_sel) begin
          accumulator_0 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_57) begin
        accumulator_1 <= io_in;
      end else begin
        accumulator_1 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h1 == io_sel) begin
          accumulator_1 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_61) begin
        accumulator_2 <= io_in;
      end else begin
        accumulator_2 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h2 == io_sel) begin
          accumulator_2 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_65) begin
        accumulator_3 <= io_in;
      end else begin
        accumulator_3 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h3 == io_sel) begin
          accumulator_3 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_69) begin
        accumulator_4 <= io_in;
      end else begin
        accumulator_4 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h4 == io_sel) begin
          accumulator_4 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_73) begin
        accumulator_5 <= io_in;
      end else begin
        accumulator_5 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h5 == io_sel) begin
          accumulator_5 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_77) begin
        accumulator_6 <= io_in;
      end else begin
        accumulator_6 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h6 == io_sel) begin
          accumulator_6 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_81) begin
        accumulator_7 <= io_in;
      end else begin
        accumulator_7 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h7 == io_sel) begin
          accumulator_7 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_85) begin
        accumulator_8 <= io_in;
      end else begin
        accumulator_8 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h8 == io_sel) begin
          accumulator_8 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_89) begin
        accumulator_9 <= io_in;
      end else begin
        accumulator_9 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h9 == io_sel) begin
          accumulator_9 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_93) begin
        accumulator_10 <= io_in;
      end else begin
        accumulator_10 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'ha == io_sel) begin
          accumulator_10 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_97) begin
        accumulator_11 <= io_in;
      end else begin
        accumulator_11 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'hb == io_sel) begin
          accumulator_11 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_101) begin
        accumulator_12 <= io_in;
      end else begin
        accumulator_12 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'hc == io_sel) begin
          accumulator_12 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_105) begin
        accumulator_13 <= io_in;
      end else begin
        accumulator_13 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'hd == io_sel) begin
          accumulator_13 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_109) begin
        accumulator_14 <= io_in;
      end else begin
        accumulator_14 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'he == io_sel) begin
          accumulator_14 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_113) begin
        accumulator_15 <= io_in;
      end else begin
        accumulator_15 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'hf == io_sel) begin
          accumulator_15 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_117) begin
        accumulator_16 <= io_in;
      end else begin
        accumulator_16 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h10 == io_sel) begin
          accumulator_16 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_121) begin
        accumulator_17 <= io_in;
      end else begin
        accumulator_17 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h11 == io_sel) begin
          accumulator_17 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_125) begin
        accumulator_18 <= io_in;
      end else begin
        accumulator_18 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h12 == io_sel) begin
          accumulator_18 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_129) begin
        accumulator_19 <= io_in;
      end else begin
        accumulator_19 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h13 == io_sel) begin
          accumulator_19 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_133) begin
        accumulator_20 <= io_in;
      end else begin
        accumulator_20 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h14 == io_sel) begin
          accumulator_20 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_137) begin
        accumulator_21 <= io_in;
      end else begin
        accumulator_21 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h15 == io_sel) begin
          accumulator_21 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_141) begin
        accumulator_22 <= io_in;
      end else begin
        accumulator_22 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h16 == io_sel) begin
          accumulator_22 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_145) begin
        accumulator_23 <= io_in;
      end else begin
        accumulator_23 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h17 == io_sel) begin
          accumulator_23 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_149) begin
        accumulator_24 <= io_in;
      end else begin
        accumulator_24 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h18 == io_sel) begin
          accumulator_24 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_153) begin
        accumulator_25 <= io_in;
      end else begin
        accumulator_25 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h19 == io_sel) begin
          accumulator_25 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_157) begin
        accumulator_26 <= io_in;
      end else begin
        accumulator_26 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h1a == io_sel) begin
          accumulator_26 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_161) begin
        accumulator_27 <= io_in;
      end else begin
        accumulator_27 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h1b == io_sel) begin
          accumulator_27 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_165) begin
        accumulator_28 <= io_in;
      end else begin
        accumulator_28 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h1c == io_sel) begin
          accumulator_28 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_169) begin
        accumulator_29 <= io_in;
      end else begin
        accumulator_29 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h1d == io_sel) begin
          accumulator_29 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_173) begin
        accumulator_30 <= io_in;
      end else begin
        accumulator_30 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h1e == io_sel) begin
          accumulator_30 <= _GEN_1;
        end
      end
    end
    if (_T_51) begin
      if (_T_177) begin
        accumulator_31 <= io_in;
      end else begin
        accumulator_31 <= 32'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h1f == io_sel) begin
          accumulator_31 <= _GEN_1;
        end
      end
    end
  end
endmodule
module MulAdd(
  input  [15:0] io_a,
  input  [15:0] io_b,
  input  [31:0] io_m,
  input  [15:0] io_c,
  output [31:0] io_r
);
  wire [31:0] _T_7;
  wire [32:0] _T_8;
  wire [32:0] _GEN_0;
  wire [64:0] _T_9;
  wire [63:0] _T_10;
  wire [63:0] _T_11;
  wire [63:0] _GEN_1;
  wire [64:0] _T_12;
  wire [63:0] _T_13;
  wire [63:0] _T_14;
  wire [31:0] _GEN_2;
  assign io_r = $signed(_GEN_2);
  assign _T_7 = $signed(io_a) * $signed(io_b);
  assign _T_8 = {1'b0,$signed(io_m)};
  assign _GEN_0 = {{1{_T_7[31]}},_T_7};
  assign _T_9 = $signed(_GEN_0) * $signed(_T_8);
  assign _T_10 = _T_9[63:0];
  assign _T_11 = $signed(_T_10);
  assign _GEN_1 = {{48{io_c[15]}},io_c};
  assign _T_12 = $signed(_T_11) + $signed(_GEN_1);
  assign _T_13 = _T_12[63:0];
  assign _T_14 = $signed(_T_13);
  assign _GEN_2 = _T_14[31:0];
endmodule
module XNORNetInference(
  input          clock,
  input          reset,
  input  [3:0]   io_input,
  input          io_inputSel,
  input          io_inputBufferPush,
  input          io_inputBufferPop,
  input          io_memSel,
  input  [7:0]   io_memAddr,
  output [127:0] io_memOut,
  input          io_memRen,
  input          io_memWen,
  input  [127:0] io_memIn,
  input          io_accEn,
  input  [4:0]   io_accSel,
  input          io_accReset,
  input          io_maxClear,
  input          io_maxEn,
  input  [3:0]   io_maxOffset,
  input          io_meanReset,
  input  [15:0]  io_featureNumInverse65536,
  input          io_meanUpdate,
  output [3:0]   io_result
);
  wire  mem_clock;
  wire [7:0] mem_io_addr;
  wire [127:0] mem_io_in;
  wire [127:0] mem_io_out;
  wire  mem_io_wen;
  wire  mem_io_ren;
  wire [3:0] inputWire;
  wire  binaryBuffer_clock;
  wire  binaryBuffer_reset;
  wire [3:0] binaryBuffer_io_in;
  wire  binaryBuffer_io_push;
  wire [31:0] binaryBuffer_io_out;
  wire  binaryBuffer_io_pop;
  wire [3:0] _T_24;
  wire [31:0] xnor$_io_in1;
  wire [31:0] xnor$_io_in2_0;
  wire [31:0] xnor$_io_in2_1;
  wire [31:0] xnor$_io_in2_2;
  wire [31:0] xnor$_io_in2_3;
  wire [31:0] xnor$_io_out_0;
  wire [31:0] xnor$_io_out_1;
  wire [31:0] xnor$_io_out_2;
  wire [31:0] xnor$_io_out_3;
  wire [31:0] _T_35_0;
  wire [31:0] _T_35_1;
  wire [31:0] _T_35_2;
  wire [31:0] _T_35_3;
  wire [127:0] _T_48;
  wire [31:0] _T_49;
  wire [31:0] _T_50;
  wire [31:0] _T_51;
  wire [31:0] _T_52;
  wire [31:0] _T_59_0;
  wire [31:0] _T_59_1;
  wire [31:0] _T_59_2;
  wire [31:0] _T_59_3;
  wire [31:0] _T_66_0;
  wire [31:0] _T_66_1;
  wire [31:0] _T_66_2;
  wire [31:0] _T_66_3;
  wire  meanBuffer_clock;
  wire  meanBuffer_reset;
  wire [31:0] meanBuffer_io_in_0;
  wire [31:0] meanBuffer_io_in_1;
  wire [31:0] meanBuffer_io_in_2;
  wire [31:0] meanBuffer_io_in_3;
  wire [15:0] meanBuffer_io_cntInverse65536;
  wire  meanBuffer_io_reset;
  wire [31:0] meanBuffer_io_out;
  wire  mean_clock;
  wire  mean_reset;
  wire [31:0] mean_io_input;
  wire  mean_io_update;
  wire [31:0] mean_io_output;
  wire  maxModule_clock;
  wire  maxModule_io_reset;
  wire  maxModule_io_en;
  wire [31:0] maxModule_io_in_0;
  wire [31:0] maxModule_io_in_1;
  wire [31:0] maxModule_io_in_2;
  wire [31:0] maxModule_io_in_3;
  wire [3:0] maxModule_io_offset;
  wire [3:0] maxModule_io_out;
  wire  Accumulator_clock;
  wire [31:0] Accumulator_io_in;
  wire [31:0] Accumulator_io_out;
  wire [4:0] Accumulator_io_sel;
  wire  Accumulator_io_en;
  wire  Accumulator_io_reset;
  wire [3:0] _T_83;
  wire [3:0] _T_84;
  wire [3:0] _T_85;
  wire [3:0] _T_86;
  wire [3:0] _T_87;
  wire [3:0] _T_88;
  wire [3:0] _T_89;
  wire [3:0] _T_90;
  reg [5:0] _T_93;
  reg [31:0] _GEN_516;
  reg [5:0] _T_96;
  reg [31:0] _GEN_517;
  reg [5:0] _T_99;
  reg [31:0] _GEN_518;
  reg [5:0] _T_102;
  reg [31:0] _GEN_519;
  reg [5:0] _T_105;
  reg [31:0] _GEN_520;
  reg [5:0] _T_108;
  reg [31:0] _GEN_521;
  reg [5:0] _T_111;
  reg [31:0] _GEN_522;
  reg [5:0] _T_114;
  reg [31:0] _GEN_523;
  reg [5:0] _T_117;
  reg [31:0] _GEN_524;
  reg [5:0] _T_120;
  reg [31:0] _GEN_525;
  reg [5:0] _T_123;
  reg [31:0] _GEN_526;
  reg [5:0] _T_126;
  reg [31:0] _GEN_527;
  reg [5:0] _T_129;
  reg [31:0] _GEN_528;
  reg [5:0] _T_132;
  reg [31:0] _GEN_529;
  reg [5:0] _T_135;
  reg [31:0] _GEN_530;
  reg [5:0] _T_138;
  reg [31:0] _GEN_531;
  wire [5:0] _T_141_0;
  wire [5:0] _T_141_1;
  wire [5:0] _T_141_2;
  wire [5:0] _T_141_3;
  wire [5:0] _T_141_4;
  wire [5:0] _T_141_5;
  wire [5:0] _T_141_6;
  wire [5:0] _T_141_7;
  wire [5:0] _T_141_8;
  wire [5:0] _T_141_9;
  wire [5:0] _T_141_10;
  wire [5:0] _T_141_11;
  wire [5:0] _T_141_12;
  wire [5:0] _T_141_13;
  wire [5:0] _T_141_14;
  wire [5:0] _T_141_15;
  reg [5:0] _T_163;
  reg [31:0] _GEN_532;
  reg [5:0] _T_166;
  reg [31:0] _GEN_533;
  reg [5:0] _T_169;
  reg [31:0] _GEN_534;
  reg [5:0] _T_172;
  reg [31:0] _GEN_535;
  reg [5:0] _T_175;
  reg [31:0] _GEN_536;
  reg [5:0] _T_178;
  reg [31:0] _GEN_537;
  reg [5:0] _T_181;
  reg [31:0] _GEN_538;
  reg [5:0] _T_184;
  reg [31:0] _GEN_539;
  reg [5:0] _T_187;
  reg [31:0] _GEN_540;
  reg [5:0] _T_190;
  reg [31:0] _GEN_541;
  reg [5:0] _T_193;
  reg [31:0] _GEN_542;
  reg [5:0] _T_196;
  reg [31:0] _GEN_543;
  reg [5:0] _T_199;
  reg [31:0] _GEN_544;
  reg [5:0] _T_202;
  reg [31:0] _GEN_545;
  reg [5:0] _T_205;
  reg [31:0] _GEN_546;
  reg [5:0] _T_208;
  reg [31:0] _GEN_547;
  wire [5:0] _T_211_0;
  wire [5:0] _T_211_1;
  wire [5:0] _T_211_2;
  wire [5:0] _T_211_3;
  wire [5:0] _T_211_4;
  wire [5:0] _T_211_5;
  wire [5:0] _T_211_6;
  wire [5:0] _T_211_7;
  wire [5:0] _T_211_8;
  wire [5:0] _T_211_9;
  wire [5:0] _T_211_10;
  wire [5:0] _T_211_11;
  wire [5:0] _T_211_12;
  wire [5:0] _T_211_13;
  wire [5:0] _T_211_14;
  wire [5:0] _T_211_15;
  reg [5:0] _T_233;
  reg [31:0] _GEN_548;
  reg [5:0] _T_236;
  reg [31:0] _GEN_549;
  reg [5:0] _T_239;
  reg [31:0] _GEN_550;
  reg [5:0] _T_242;
  reg [31:0] _GEN_551;
  reg [5:0] _T_245;
  reg [31:0] _GEN_552;
  reg [5:0] _T_248;
  reg [31:0] _GEN_553;
  reg [5:0] _T_251;
  reg [31:0] _GEN_554;
  reg [5:0] _T_254;
  reg [31:0] _GEN_555;
  reg [5:0] _T_257;
  reg [31:0] _GEN_556;
  reg [5:0] _T_260;
  reg [31:0] _GEN_557;
  reg [5:0] _T_263;
  reg [31:0] _GEN_558;
  reg [5:0] _T_266;
  reg [31:0] _GEN_559;
  reg [5:0] _T_269;
  reg [31:0] _GEN_560;
  reg [5:0] _T_272;
  reg [31:0] _GEN_561;
  reg [5:0] _T_275;
  reg [31:0] _GEN_562;
  reg [5:0] _T_278;
  reg [31:0] _GEN_563;
  wire [5:0] _T_281_0;
  wire [5:0] _T_281_1;
  wire [5:0] _T_281_2;
  wire [5:0] _T_281_3;
  wire [5:0] _T_281_4;
  wire [5:0] _T_281_5;
  wire [5:0] _T_281_6;
  wire [5:0] _T_281_7;
  wire [5:0] _T_281_8;
  wire [5:0] _T_281_9;
  wire [5:0] _T_281_10;
  wire [5:0] _T_281_11;
  wire [5:0] _T_281_12;
  wire [5:0] _T_281_13;
  wire [5:0] _T_281_14;
  wire [5:0] _T_281_15;
  reg [5:0] _T_303;
  reg [31:0] _GEN_564;
  reg [5:0] _T_306;
  reg [31:0] _GEN_565;
  reg [5:0] _T_309;
  reg [31:0] _GEN_566;
  reg [5:0] _T_312;
  reg [31:0] _GEN_567;
  reg [5:0] _T_315;
  reg [31:0] _GEN_568;
  reg [5:0] _T_318;
  reg [31:0] _GEN_569;
  reg [5:0] _T_321;
  reg [31:0] _GEN_570;
  reg [5:0] _T_324;
  reg [31:0] _GEN_571;
  reg [5:0] _T_327;
  reg [31:0] _GEN_572;
  reg [5:0] _T_330;
  reg [31:0] _GEN_573;
  reg [5:0] _T_333;
  reg [31:0] _GEN_574;
  reg [5:0] _T_336;
  reg [31:0] _GEN_575;
  reg [5:0] _T_339;
  reg [31:0] _GEN_576;
  reg [5:0] _T_342;
  reg [31:0] _GEN_577;
  reg [5:0] _T_345;
  reg [31:0] _GEN_578;
  reg [5:0] _T_348;
  reg [31:0] _GEN_579;
  wire [5:0] _T_351_0;
  wire [5:0] _T_351_1;
  wire [5:0] _T_351_2;
  wire [5:0] _T_351_3;
  wire [5:0] _T_351_4;
  wire [5:0] _T_351_5;
  wire [5:0] _T_351_6;
  wire [5:0] _T_351_7;
  wire [5:0] _T_351_8;
  wire [5:0] _T_351_9;
  wire [5:0] _T_351_10;
  wire [5:0] _T_351_11;
  wire [5:0] _T_351_12;
  wire [5:0] _T_351_13;
  wire [5:0] _T_351_14;
  wire [5:0] _T_351_15;
  reg [5:0] _T_373;
  reg [31:0] _GEN_580;
  reg [5:0] _T_376;
  reg [31:0] _GEN_581;
  reg [5:0] _T_379;
  reg [31:0] _GEN_582;
  reg [5:0] _T_382;
  reg [31:0] _GEN_583;
  reg [5:0] _T_385;
  reg [31:0] _GEN_584;
  reg [5:0] _T_388;
  reg [31:0] _GEN_585;
  reg [5:0] _T_391;
  reg [31:0] _GEN_586;
  reg [5:0] _T_394;
  reg [31:0] _GEN_587;
  reg [5:0] _T_397;
  reg [31:0] _GEN_588;
  reg [5:0] _T_400;
  reg [31:0] _GEN_589;
  reg [5:0] _T_403;
  reg [31:0] _GEN_590;
  reg [5:0] _T_406;
  reg [31:0] _GEN_591;
  reg [5:0] _T_409;
  reg [31:0] _GEN_592;
  reg [5:0] _T_412;
  reg [31:0] _GEN_593;
  reg [5:0] _T_415;
  reg [31:0] _GEN_594;
  reg [5:0] _T_418;
  reg [31:0] _GEN_595;
  wire [5:0] _T_421_0;
  wire [5:0] _T_421_1;
  wire [5:0] _T_421_2;
  wire [5:0] _T_421_3;
  wire [5:0] _T_421_4;
  wire [5:0] _T_421_5;
  wire [5:0] _T_421_6;
  wire [5:0] _T_421_7;
  wire [5:0] _T_421_8;
  wire [5:0] _T_421_9;
  wire [5:0] _T_421_10;
  wire [5:0] _T_421_11;
  wire [5:0] _T_421_12;
  wire [5:0] _T_421_13;
  wire [5:0] _T_421_14;
  wire [5:0] _T_421_15;
  reg [5:0] _T_443;
  reg [31:0] _GEN_596;
  reg [5:0] _T_446;
  reg [31:0] _GEN_597;
  reg [5:0] _T_449;
  reg [31:0] _GEN_598;
  reg [5:0] _T_452;
  reg [31:0] _GEN_599;
  reg [5:0] _T_455;
  reg [31:0] _GEN_600;
  reg [5:0] _T_458;
  reg [31:0] _GEN_601;
  reg [5:0] _T_461;
  reg [31:0] _GEN_602;
  reg [5:0] _T_464;
  reg [31:0] _GEN_603;
  reg [5:0] _T_467;
  reg [31:0] _GEN_604;
  reg [5:0] _T_470;
  reg [31:0] _GEN_605;
  reg [5:0] _T_473;
  reg [31:0] _GEN_606;
  reg [5:0] _T_476;
  reg [31:0] _GEN_607;
  reg [5:0] _T_479;
  reg [31:0] _GEN_608;
  reg [5:0] _T_482;
  reg [31:0] _GEN_609;
  reg [5:0] _T_485;
  reg [31:0] _GEN_610;
  reg [5:0] _T_488;
  reg [31:0] _GEN_611;
  wire [5:0] _T_491_0;
  wire [5:0] _T_491_1;
  wire [5:0] _T_491_2;
  wire [5:0] _T_491_3;
  wire [5:0] _T_491_4;
  wire [5:0] _T_491_5;
  wire [5:0] _T_491_6;
  wire [5:0] _T_491_7;
  wire [5:0] _T_491_8;
  wire [5:0] _T_491_9;
  wire [5:0] _T_491_10;
  wire [5:0] _T_491_11;
  wire [5:0] _T_491_12;
  wire [5:0] _T_491_13;
  wire [5:0] _T_491_14;
  wire [5:0] _T_491_15;
  reg [5:0] _T_513;
  reg [31:0] _GEN_612;
  reg [5:0] _T_516;
  reg [31:0] _GEN_613;
  reg [5:0] _T_519;
  reg [31:0] _GEN_614;
  reg [5:0] _T_522;
  reg [31:0] _GEN_615;
  reg [5:0] _T_525;
  reg [31:0] _GEN_616;
  reg [5:0] _T_528;
  reg [31:0] _GEN_617;
  reg [5:0] _T_531;
  reg [31:0] _GEN_618;
  reg [5:0] _T_534;
  reg [31:0] _GEN_619;
  reg [5:0] _T_537;
  reg [31:0] _GEN_620;
  reg [5:0] _T_540;
  reg [31:0] _GEN_621;
  reg [5:0] _T_543;
  reg [31:0] _GEN_622;
  reg [5:0] _T_546;
  reg [31:0] _GEN_623;
  reg [5:0] _T_549;
  reg [31:0] _GEN_624;
  reg [5:0] _T_552;
  reg [31:0] _GEN_625;
  reg [5:0] _T_555;
  reg [31:0] _GEN_626;
  reg [5:0] _T_558;
  reg [31:0] _GEN_627;
  wire [5:0] _T_561_0;
  wire [5:0] _T_561_1;
  wire [5:0] _T_561_2;
  wire [5:0] _T_561_3;
  wire [5:0] _T_561_4;
  wire [5:0] _T_561_5;
  wire [5:0] _T_561_6;
  wire [5:0] _T_561_7;
  wire [5:0] _T_561_8;
  wire [5:0] _T_561_9;
  wire [5:0] _T_561_10;
  wire [5:0] _T_561_11;
  wire [5:0] _T_561_12;
  wire [5:0] _T_561_13;
  wire [5:0] _T_561_14;
  wire [5:0] _T_561_15;
  reg [5:0] _T_583;
  reg [31:0] _GEN_628;
  reg [5:0] _T_586;
  reg [31:0] _GEN_629;
  reg [5:0] _T_589;
  reg [31:0] _GEN_630;
  reg [5:0] _T_592;
  reg [31:0] _GEN_631;
  reg [5:0] _T_595;
  reg [31:0] _GEN_632;
  reg [5:0] _T_598;
  reg [31:0] _GEN_633;
  reg [5:0] _T_601;
  reg [31:0] _GEN_634;
  reg [5:0] _T_604;
  reg [31:0] _GEN_635;
  reg [5:0] _T_607;
  reg [31:0] _GEN_636;
  reg [5:0] _T_610;
  reg [31:0] _GEN_637;
  reg [5:0] _T_613;
  reg [31:0] _GEN_638;
  reg [5:0] _T_616;
  reg [31:0] _GEN_639;
  reg [5:0] _T_619;
  reg [31:0] _GEN_640;
  reg [5:0] _T_622;
  reg [31:0] _GEN_641;
  reg [5:0] _T_625;
  reg [31:0] _GEN_642;
  reg [5:0] _T_628;
  reg [31:0] _GEN_643;
  wire [5:0] _T_631_0;
  wire [5:0] _T_631_1;
  wire [5:0] _T_631_2;
  wire [5:0] _T_631_3;
  wire [5:0] _T_631_4;
  wire [5:0] _T_631_5;
  wire [5:0] _T_631_6;
  wire [5:0] _T_631_7;
  wire [5:0] _T_631_8;
  wire [5:0] _T_631_9;
  wire [5:0] _T_631_10;
  wire [5:0] _T_631_11;
  wire [5:0] _T_631_12;
  wire [5:0] _T_631_13;
  wire [5:0] _T_631_14;
  wire [5:0] _T_631_15;
  wire [5:0] _GEN_0;
  wire [5:0] _GEN_32;
  wire [5:0] _GEN_33;
  wire [5:0] _GEN_34;
  wire [5:0] _GEN_35;
  wire [5:0] _GEN_36;
  wire [5:0] _GEN_37;
  wire [5:0] _GEN_38;
  wire [5:0] _GEN_39;
  wire [5:0] _GEN_40;
  wire [5:0] _GEN_41;
  wire [5:0] _GEN_42;
  wire [5:0] _GEN_43;
  wire [5:0] _GEN_44;
  wire [5:0] _GEN_45;
  wire [5:0] _GEN_46;
  wire [5:0] _GEN_1;
  wire [5:0] _GEN_47;
  wire [5:0] _GEN_48;
  wire [5:0] _GEN_49;
  wire [5:0] _GEN_50;
  wire [5:0] _GEN_51;
  wire [5:0] _GEN_52;
  wire [5:0] _GEN_53;
  wire [5:0] _GEN_54;
  wire [5:0] _GEN_55;
  wire [5:0] _GEN_56;
  wire [5:0] _GEN_57;
  wire [5:0] _GEN_58;
  wire [5:0] _GEN_59;
  wire [5:0] _GEN_60;
  wire [5:0] _GEN_61;
  wire [6:0] _T_651;
  wire [5:0] _T_652;
  wire [5:0] _T_653;
  wire [5:0] _GEN_2;
  wire [5:0] _GEN_62;
  wire [5:0] _GEN_63;
  wire [5:0] _GEN_64;
  wire [5:0] _GEN_65;
  wire [5:0] _GEN_66;
  wire [5:0] _GEN_67;
  wire [5:0] _GEN_68;
  wire [5:0] _GEN_69;
  wire [5:0] _GEN_70;
  wire [5:0] _GEN_71;
  wire [5:0] _GEN_72;
  wire [5:0] _GEN_73;
  wire [5:0] _GEN_74;
  wire [5:0] _GEN_75;
  wire [5:0] _GEN_76;
  wire [5:0] _GEN_3;
  wire [5:0] _GEN_77;
  wire [5:0] _GEN_78;
  wire [5:0] _GEN_79;
  wire [5:0] _GEN_80;
  wire [5:0] _GEN_81;
  wire [5:0] _GEN_82;
  wire [5:0] _GEN_83;
  wire [5:0] _GEN_84;
  wire [5:0] _GEN_85;
  wire [5:0] _GEN_86;
  wire [5:0] _GEN_87;
  wire [5:0] _GEN_88;
  wire [5:0] _GEN_89;
  wire [5:0] _GEN_90;
  wire [5:0] _GEN_91;
  wire [6:0] _T_654;
  wire [5:0] _T_655;
  wire [5:0] _T_656;
  wire [5:0] _GEN_4;
  wire [5:0] _GEN_92;
  wire [5:0] _GEN_93;
  wire [5:0] _GEN_94;
  wire [5:0] _GEN_95;
  wire [5:0] _GEN_96;
  wire [5:0] _GEN_97;
  wire [5:0] _GEN_98;
  wire [5:0] _GEN_99;
  wire [5:0] _GEN_100;
  wire [5:0] _GEN_101;
  wire [5:0] _GEN_102;
  wire [5:0] _GEN_103;
  wire [5:0] _GEN_104;
  wire [5:0] _GEN_105;
  wire [5:0] _GEN_106;
  wire [5:0] _GEN_5;
  wire [5:0] _GEN_107;
  wire [5:0] _GEN_108;
  wire [5:0] _GEN_109;
  wire [5:0] _GEN_110;
  wire [5:0] _GEN_111;
  wire [5:0] _GEN_112;
  wire [5:0] _GEN_113;
  wire [5:0] _GEN_114;
  wire [5:0] _GEN_115;
  wire [5:0] _GEN_116;
  wire [5:0] _GEN_117;
  wire [5:0] _GEN_118;
  wire [5:0] _GEN_119;
  wire [5:0] _GEN_120;
  wire [5:0] _GEN_121;
  wire [6:0] _T_657;
  wire [5:0] _T_658;
  wire [5:0] _T_659;
  wire [5:0] _GEN_6;
  wire [5:0] _GEN_122;
  wire [5:0] _GEN_123;
  wire [5:0] _GEN_124;
  wire [5:0] _GEN_125;
  wire [5:0] _GEN_126;
  wire [5:0] _GEN_127;
  wire [5:0] _GEN_128;
  wire [5:0] _GEN_129;
  wire [5:0] _GEN_130;
  wire [5:0] _GEN_131;
  wire [5:0] _GEN_132;
  wire [5:0] _GEN_133;
  wire [5:0] _GEN_134;
  wire [5:0] _GEN_135;
  wire [5:0] _GEN_136;
  wire [5:0] _GEN_7;
  wire [5:0] _GEN_137;
  wire [5:0] _GEN_138;
  wire [5:0] _GEN_139;
  wire [5:0] _GEN_140;
  wire [5:0] _GEN_141;
  wire [5:0] _GEN_142;
  wire [5:0] _GEN_143;
  wire [5:0] _GEN_144;
  wire [5:0] _GEN_145;
  wire [5:0] _GEN_146;
  wire [5:0] _GEN_147;
  wire [5:0] _GEN_148;
  wire [5:0] _GEN_149;
  wire [5:0] _GEN_150;
  wire [5:0] _GEN_151;
  wire [6:0] _T_660;
  wire [5:0] _T_661;
  wire [5:0] _T_662;
  wire [6:0] _T_663;
  wire [5:0] _T_664;
  wire [5:0] _T_665;
  wire [6:0] _T_666;
  wire [5:0] _T_667;
  wire [5:0] _T_668;
  wire [6:0] _T_669;
  wire [5:0] _T_670;
  wire [5:0] _T_671;
  wire [15:0] MulAdd_io_a;
  wire [15:0] MulAdd_io_b;
  wire [31:0] MulAdd_io_m;
  wire [15:0] MulAdd_io_c;
  wire [31:0] MulAdd_io_r;
  wire [31:0] _T_673;
  wire [31:0] _T_674;
  wire [15:0] _T_675;
  wire [15:0] _T_676;
  wire [15:0] _T_677;
  wire [15:0] _T_678;
  wire  signs_0;
  wire  Accumulator_1_clock;
  wire [31:0] Accumulator_1_io_in;
  wire [31:0] Accumulator_1_io_out;
  wire [4:0] Accumulator_1_io_sel;
  wire  Accumulator_1_io_en;
  wire  Accumulator_1_io_reset;
  wire [3:0] _T_679;
  wire [3:0] _T_680;
  wire [3:0] _T_681;
  wire [3:0] _T_682;
  wire [3:0] _T_683;
  wire [3:0] _T_684;
  wire [3:0] _T_685;
  wire [3:0] _T_686;
  reg [5:0] _T_689;
  reg [31:0] _GEN_644;
  reg [5:0] _T_692;
  reg [31:0] _GEN_645;
  reg [5:0] _T_695;
  reg [31:0] _GEN_646;
  reg [5:0] _T_698;
  reg [31:0] _GEN_647;
  reg [5:0] _T_701;
  reg [31:0] _GEN_648;
  reg [5:0] _T_704;
  reg [31:0] _GEN_649;
  reg [5:0] _T_707;
  reg [31:0] _GEN_650;
  reg [5:0] _T_710;
  reg [31:0] _GEN_651;
  reg [5:0] _T_713;
  reg [31:0] _GEN_652;
  reg [5:0] _T_716;
  reg [31:0] _GEN_653;
  reg [5:0] _T_719;
  reg [31:0] _GEN_654;
  reg [5:0] _T_722;
  reg [31:0] _GEN_655;
  reg [5:0] _T_725;
  reg [31:0] _GEN_656;
  reg [5:0] _T_728;
  reg [31:0] _GEN_657;
  reg [5:0] _T_731;
  reg [31:0] _GEN_658;
  reg [5:0] _T_734;
  reg [31:0] _GEN_659;
  wire [5:0] _T_737_0;
  wire [5:0] _T_737_1;
  wire [5:0] _T_737_2;
  wire [5:0] _T_737_3;
  wire [5:0] _T_737_4;
  wire [5:0] _T_737_5;
  wire [5:0] _T_737_6;
  wire [5:0] _T_737_7;
  wire [5:0] _T_737_8;
  wire [5:0] _T_737_9;
  wire [5:0] _T_737_10;
  wire [5:0] _T_737_11;
  wire [5:0] _T_737_12;
  wire [5:0] _T_737_13;
  wire [5:0] _T_737_14;
  wire [5:0] _T_737_15;
  reg [5:0] _T_759;
  reg [31:0] _GEN_660;
  reg [5:0] _T_762;
  reg [31:0] _GEN_661;
  reg [5:0] _T_765;
  reg [31:0] _GEN_662;
  reg [5:0] _T_768;
  reg [31:0] _GEN_663;
  reg [5:0] _T_771;
  reg [31:0] _GEN_664;
  reg [5:0] _T_774;
  reg [31:0] _GEN_665;
  reg [5:0] _T_777;
  reg [31:0] _GEN_666;
  reg [5:0] _T_780;
  reg [31:0] _GEN_667;
  reg [5:0] _T_783;
  reg [31:0] _GEN_668;
  reg [5:0] _T_786;
  reg [31:0] _GEN_669;
  reg [5:0] _T_789;
  reg [31:0] _GEN_670;
  reg [5:0] _T_792;
  reg [31:0] _GEN_671;
  reg [5:0] _T_795;
  reg [31:0] _GEN_672;
  reg [5:0] _T_798;
  reg [31:0] _GEN_673;
  reg [5:0] _T_801;
  reg [31:0] _GEN_674;
  reg [5:0] _T_804;
  reg [31:0] _GEN_675;
  wire [5:0] _T_807_0;
  wire [5:0] _T_807_1;
  wire [5:0] _T_807_2;
  wire [5:0] _T_807_3;
  wire [5:0] _T_807_4;
  wire [5:0] _T_807_5;
  wire [5:0] _T_807_6;
  wire [5:0] _T_807_7;
  wire [5:0] _T_807_8;
  wire [5:0] _T_807_9;
  wire [5:0] _T_807_10;
  wire [5:0] _T_807_11;
  wire [5:0] _T_807_12;
  wire [5:0] _T_807_13;
  wire [5:0] _T_807_14;
  wire [5:0] _T_807_15;
  reg [5:0] _T_829;
  reg [31:0] _GEN_676;
  reg [5:0] _T_832;
  reg [31:0] _GEN_677;
  reg [5:0] _T_835;
  reg [31:0] _GEN_678;
  reg [5:0] _T_838;
  reg [31:0] _GEN_679;
  reg [5:0] _T_841;
  reg [31:0] _GEN_680;
  reg [5:0] _T_844;
  reg [31:0] _GEN_681;
  reg [5:0] _T_847;
  reg [31:0] _GEN_682;
  reg [5:0] _T_850;
  reg [31:0] _GEN_683;
  reg [5:0] _T_853;
  reg [31:0] _GEN_684;
  reg [5:0] _T_856;
  reg [31:0] _GEN_685;
  reg [5:0] _T_859;
  reg [31:0] _GEN_686;
  reg [5:0] _T_862;
  reg [31:0] _GEN_687;
  reg [5:0] _T_865;
  reg [31:0] _GEN_688;
  reg [5:0] _T_868;
  reg [31:0] _GEN_689;
  reg [5:0] _T_871;
  reg [31:0] _GEN_690;
  reg [5:0] _T_874;
  reg [31:0] _GEN_691;
  wire [5:0] _T_877_0;
  wire [5:0] _T_877_1;
  wire [5:0] _T_877_2;
  wire [5:0] _T_877_3;
  wire [5:0] _T_877_4;
  wire [5:0] _T_877_5;
  wire [5:0] _T_877_6;
  wire [5:0] _T_877_7;
  wire [5:0] _T_877_8;
  wire [5:0] _T_877_9;
  wire [5:0] _T_877_10;
  wire [5:0] _T_877_11;
  wire [5:0] _T_877_12;
  wire [5:0] _T_877_13;
  wire [5:0] _T_877_14;
  wire [5:0] _T_877_15;
  reg [5:0] _T_899;
  reg [31:0] _GEN_692;
  reg [5:0] _T_902;
  reg [31:0] _GEN_693;
  reg [5:0] _T_905;
  reg [31:0] _GEN_694;
  reg [5:0] _T_908;
  reg [31:0] _GEN_695;
  reg [5:0] _T_911;
  reg [31:0] _GEN_696;
  reg [5:0] _T_914;
  reg [31:0] _GEN_697;
  reg [5:0] _T_917;
  reg [31:0] _GEN_698;
  reg [5:0] _T_920;
  reg [31:0] _GEN_699;
  reg [5:0] _T_923;
  reg [31:0] _GEN_700;
  reg [5:0] _T_926;
  reg [31:0] _GEN_701;
  reg [5:0] _T_929;
  reg [31:0] _GEN_702;
  reg [5:0] _T_932;
  reg [31:0] _GEN_703;
  reg [5:0] _T_935;
  reg [31:0] _GEN_704;
  reg [5:0] _T_938;
  reg [31:0] _GEN_705;
  reg [5:0] _T_941;
  reg [31:0] _GEN_706;
  reg [5:0] _T_944;
  reg [31:0] _GEN_707;
  wire [5:0] _T_947_0;
  wire [5:0] _T_947_1;
  wire [5:0] _T_947_2;
  wire [5:0] _T_947_3;
  wire [5:0] _T_947_4;
  wire [5:0] _T_947_5;
  wire [5:0] _T_947_6;
  wire [5:0] _T_947_7;
  wire [5:0] _T_947_8;
  wire [5:0] _T_947_9;
  wire [5:0] _T_947_10;
  wire [5:0] _T_947_11;
  wire [5:0] _T_947_12;
  wire [5:0] _T_947_13;
  wire [5:0] _T_947_14;
  wire [5:0] _T_947_15;
  reg [5:0] _T_969;
  reg [31:0] _GEN_708;
  reg [5:0] _T_972;
  reg [31:0] _GEN_709;
  reg [5:0] _T_975;
  reg [31:0] _GEN_710;
  reg [5:0] _T_978;
  reg [31:0] _GEN_711;
  reg [5:0] _T_981;
  reg [31:0] _GEN_712;
  reg [5:0] _T_984;
  reg [31:0] _GEN_713;
  reg [5:0] _T_987;
  reg [31:0] _GEN_714;
  reg [5:0] _T_990;
  reg [31:0] _GEN_715;
  reg [5:0] _T_993;
  reg [31:0] _GEN_716;
  reg [5:0] _T_996;
  reg [31:0] _GEN_717;
  reg [5:0] _T_999;
  reg [31:0] _GEN_718;
  reg [5:0] _T_1002;
  reg [31:0] _GEN_719;
  reg [5:0] _T_1005;
  reg [31:0] _GEN_720;
  reg [5:0] _T_1008;
  reg [31:0] _GEN_721;
  reg [5:0] _T_1011;
  reg [31:0] _GEN_722;
  reg [5:0] _T_1014;
  reg [31:0] _GEN_723;
  wire [5:0] _T_1017_0;
  wire [5:0] _T_1017_1;
  wire [5:0] _T_1017_2;
  wire [5:0] _T_1017_3;
  wire [5:0] _T_1017_4;
  wire [5:0] _T_1017_5;
  wire [5:0] _T_1017_6;
  wire [5:0] _T_1017_7;
  wire [5:0] _T_1017_8;
  wire [5:0] _T_1017_9;
  wire [5:0] _T_1017_10;
  wire [5:0] _T_1017_11;
  wire [5:0] _T_1017_12;
  wire [5:0] _T_1017_13;
  wire [5:0] _T_1017_14;
  wire [5:0] _T_1017_15;
  reg [5:0] _T_1039;
  reg [31:0] _GEN_724;
  reg [5:0] _T_1042;
  reg [31:0] _GEN_725;
  reg [5:0] _T_1045;
  reg [31:0] _GEN_726;
  reg [5:0] _T_1048;
  reg [31:0] _GEN_727;
  reg [5:0] _T_1051;
  reg [31:0] _GEN_728;
  reg [5:0] _T_1054;
  reg [31:0] _GEN_729;
  reg [5:0] _T_1057;
  reg [31:0] _GEN_730;
  reg [5:0] _T_1060;
  reg [31:0] _GEN_731;
  reg [5:0] _T_1063;
  reg [31:0] _GEN_732;
  reg [5:0] _T_1066;
  reg [31:0] _GEN_733;
  reg [5:0] _T_1069;
  reg [31:0] _GEN_734;
  reg [5:0] _T_1072;
  reg [31:0] _GEN_735;
  reg [5:0] _T_1075;
  reg [31:0] _GEN_736;
  reg [5:0] _T_1078;
  reg [31:0] _GEN_737;
  reg [5:0] _T_1081;
  reg [31:0] _GEN_738;
  reg [5:0] _T_1084;
  reg [31:0] _GEN_739;
  wire [5:0] _T_1087_0;
  wire [5:0] _T_1087_1;
  wire [5:0] _T_1087_2;
  wire [5:0] _T_1087_3;
  wire [5:0] _T_1087_4;
  wire [5:0] _T_1087_5;
  wire [5:0] _T_1087_6;
  wire [5:0] _T_1087_7;
  wire [5:0] _T_1087_8;
  wire [5:0] _T_1087_9;
  wire [5:0] _T_1087_10;
  wire [5:0] _T_1087_11;
  wire [5:0] _T_1087_12;
  wire [5:0] _T_1087_13;
  wire [5:0] _T_1087_14;
  wire [5:0] _T_1087_15;
  reg [5:0] _T_1109;
  reg [31:0] _GEN_740;
  reg [5:0] _T_1112;
  reg [31:0] _GEN_741;
  reg [5:0] _T_1115;
  reg [31:0] _GEN_742;
  reg [5:0] _T_1118;
  reg [31:0] _GEN_743;
  reg [5:0] _T_1121;
  reg [31:0] _GEN_744;
  reg [5:0] _T_1124;
  reg [31:0] _GEN_745;
  reg [5:0] _T_1127;
  reg [31:0] _GEN_746;
  reg [5:0] _T_1130;
  reg [31:0] _GEN_747;
  reg [5:0] _T_1133;
  reg [31:0] _GEN_748;
  reg [5:0] _T_1136;
  reg [31:0] _GEN_749;
  reg [5:0] _T_1139;
  reg [31:0] _GEN_750;
  reg [5:0] _T_1142;
  reg [31:0] _GEN_751;
  reg [5:0] _T_1145;
  reg [31:0] _GEN_752;
  reg [5:0] _T_1148;
  reg [31:0] _GEN_753;
  reg [5:0] _T_1151;
  reg [31:0] _GEN_754;
  reg [5:0] _T_1154;
  reg [31:0] _GEN_755;
  wire [5:0] _T_1157_0;
  wire [5:0] _T_1157_1;
  wire [5:0] _T_1157_2;
  wire [5:0] _T_1157_3;
  wire [5:0] _T_1157_4;
  wire [5:0] _T_1157_5;
  wire [5:0] _T_1157_6;
  wire [5:0] _T_1157_7;
  wire [5:0] _T_1157_8;
  wire [5:0] _T_1157_9;
  wire [5:0] _T_1157_10;
  wire [5:0] _T_1157_11;
  wire [5:0] _T_1157_12;
  wire [5:0] _T_1157_13;
  wire [5:0] _T_1157_14;
  wire [5:0] _T_1157_15;
  reg [5:0] _T_1179;
  reg [31:0] _GEN_756;
  reg [5:0] _T_1182;
  reg [31:0] _GEN_757;
  reg [5:0] _T_1185;
  reg [31:0] _GEN_758;
  reg [5:0] _T_1188;
  reg [31:0] _GEN_759;
  reg [5:0] _T_1191;
  reg [31:0] _GEN_760;
  reg [5:0] _T_1194;
  reg [31:0] _GEN_761;
  reg [5:0] _T_1197;
  reg [31:0] _GEN_762;
  reg [5:0] _T_1200;
  reg [31:0] _GEN_763;
  reg [5:0] _T_1203;
  reg [31:0] _GEN_764;
  reg [5:0] _T_1206;
  reg [31:0] _GEN_765;
  reg [5:0] _T_1209;
  reg [31:0] _GEN_766;
  reg [5:0] _T_1212;
  reg [31:0] _GEN_767;
  reg [5:0] _T_1215;
  reg [31:0] _GEN_768;
  reg [5:0] _T_1218;
  reg [31:0] _GEN_769;
  reg [5:0] _T_1221;
  reg [31:0] _GEN_770;
  reg [5:0] _T_1224;
  reg [31:0] _GEN_771;
  wire [5:0] _T_1227_0;
  wire [5:0] _T_1227_1;
  wire [5:0] _T_1227_2;
  wire [5:0] _T_1227_3;
  wire [5:0] _T_1227_4;
  wire [5:0] _T_1227_5;
  wire [5:0] _T_1227_6;
  wire [5:0] _T_1227_7;
  wire [5:0] _T_1227_8;
  wire [5:0] _T_1227_9;
  wire [5:0] _T_1227_10;
  wire [5:0] _T_1227_11;
  wire [5:0] _T_1227_12;
  wire [5:0] _T_1227_13;
  wire [5:0] _T_1227_14;
  wire [5:0] _T_1227_15;
  wire [5:0] _GEN_8;
  wire [5:0] _GEN_152;
  wire [5:0] _GEN_153;
  wire [5:0] _GEN_154;
  wire [5:0] _GEN_155;
  wire [5:0] _GEN_156;
  wire [5:0] _GEN_157;
  wire [5:0] _GEN_158;
  wire [5:0] _GEN_159;
  wire [5:0] _GEN_160;
  wire [5:0] _GEN_161;
  wire [5:0] _GEN_162;
  wire [5:0] _GEN_163;
  wire [5:0] _GEN_164;
  wire [5:0] _GEN_165;
  wire [5:0] _GEN_166;
  wire [5:0] _GEN_9;
  wire [5:0] _GEN_167;
  wire [5:0] _GEN_168;
  wire [5:0] _GEN_169;
  wire [5:0] _GEN_170;
  wire [5:0] _GEN_171;
  wire [5:0] _GEN_172;
  wire [5:0] _GEN_173;
  wire [5:0] _GEN_174;
  wire [5:0] _GEN_175;
  wire [5:0] _GEN_176;
  wire [5:0] _GEN_177;
  wire [5:0] _GEN_178;
  wire [5:0] _GEN_179;
  wire [5:0] _GEN_180;
  wire [5:0] _GEN_181;
  wire [6:0] _T_1247;
  wire [5:0] _T_1248;
  wire [5:0] _T_1249;
  wire [5:0] _GEN_10;
  wire [5:0] _GEN_182;
  wire [5:0] _GEN_183;
  wire [5:0] _GEN_184;
  wire [5:0] _GEN_185;
  wire [5:0] _GEN_186;
  wire [5:0] _GEN_187;
  wire [5:0] _GEN_188;
  wire [5:0] _GEN_189;
  wire [5:0] _GEN_190;
  wire [5:0] _GEN_191;
  wire [5:0] _GEN_192;
  wire [5:0] _GEN_193;
  wire [5:0] _GEN_194;
  wire [5:0] _GEN_195;
  wire [5:0] _GEN_196;
  wire [5:0] _GEN_11;
  wire [5:0] _GEN_197;
  wire [5:0] _GEN_198;
  wire [5:0] _GEN_199;
  wire [5:0] _GEN_200;
  wire [5:0] _GEN_201;
  wire [5:0] _GEN_202;
  wire [5:0] _GEN_203;
  wire [5:0] _GEN_204;
  wire [5:0] _GEN_205;
  wire [5:0] _GEN_206;
  wire [5:0] _GEN_207;
  wire [5:0] _GEN_208;
  wire [5:0] _GEN_209;
  wire [5:0] _GEN_210;
  wire [5:0] _GEN_211;
  wire [6:0] _T_1250;
  wire [5:0] _T_1251;
  wire [5:0] _T_1252;
  wire [5:0] _GEN_12;
  wire [5:0] _GEN_212;
  wire [5:0] _GEN_213;
  wire [5:0] _GEN_214;
  wire [5:0] _GEN_215;
  wire [5:0] _GEN_216;
  wire [5:0] _GEN_217;
  wire [5:0] _GEN_218;
  wire [5:0] _GEN_219;
  wire [5:0] _GEN_220;
  wire [5:0] _GEN_221;
  wire [5:0] _GEN_222;
  wire [5:0] _GEN_223;
  wire [5:0] _GEN_224;
  wire [5:0] _GEN_225;
  wire [5:0] _GEN_226;
  wire [5:0] _GEN_13;
  wire [5:0] _GEN_227;
  wire [5:0] _GEN_228;
  wire [5:0] _GEN_229;
  wire [5:0] _GEN_230;
  wire [5:0] _GEN_231;
  wire [5:0] _GEN_232;
  wire [5:0] _GEN_233;
  wire [5:0] _GEN_234;
  wire [5:0] _GEN_235;
  wire [5:0] _GEN_236;
  wire [5:0] _GEN_237;
  wire [5:0] _GEN_238;
  wire [5:0] _GEN_239;
  wire [5:0] _GEN_240;
  wire [5:0] _GEN_241;
  wire [6:0] _T_1253;
  wire [5:0] _T_1254;
  wire [5:0] _T_1255;
  wire [5:0] _GEN_14;
  wire [5:0] _GEN_242;
  wire [5:0] _GEN_243;
  wire [5:0] _GEN_244;
  wire [5:0] _GEN_245;
  wire [5:0] _GEN_246;
  wire [5:0] _GEN_247;
  wire [5:0] _GEN_248;
  wire [5:0] _GEN_249;
  wire [5:0] _GEN_250;
  wire [5:0] _GEN_251;
  wire [5:0] _GEN_252;
  wire [5:0] _GEN_253;
  wire [5:0] _GEN_254;
  wire [5:0] _GEN_255;
  wire [5:0] _GEN_256;
  wire [5:0] _GEN_15;
  wire [5:0] _GEN_257;
  wire [5:0] _GEN_258;
  wire [5:0] _GEN_259;
  wire [5:0] _GEN_260;
  wire [5:0] _GEN_261;
  wire [5:0] _GEN_262;
  wire [5:0] _GEN_263;
  wire [5:0] _GEN_264;
  wire [5:0] _GEN_265;
  wire [5:0] _GEN_266;
  wire [5:0] _GEN_267;
  wire [5:0] _GEN_268;
  wire [5:0] _GEN_269;
  wire [5:0] _GEN_270;
  wire [5:0] _GEN_271;
  wire [6:0] _T_1256;
  wire [5:0] _T_1257;
  wire [5:0] _T_1258;
  wire [6:0] _T_1259;
  wire [5:0] _T_1260;
  wire [5:0] _T_1261;
  wire [6:0] _T_1262;
  wire [5:0] _T_1263;
  wire [5:0] _T_1264;
  wire [6:0] _T_1265;
  wire [5:0] _T_1266;
  wire [5:0] _T_1267;
  wire [15:0] MulAdd_1_io_a;
  wire [15:0] MulAdd_1_io_b;
  wire [31:0] MulAdd_1_io_m;
  wire [15:0] MulAdd_1_io_c;
  wire [31:0] MulAdd_1_io_r;
  wire [31:0] _T_1269;
  wire [31:0] _T_1270;
  wire [15:0] _T_1271;
  wire [15:0] _T_1272;
  wire [15:0] _T_1273;
  wire [15:0] _T_1274;
  wire  signs_1;
  wire  Accumulator_2_clock;
  wire [31:0] Accumulator_2_io_in;
  wire [31:0] Accumulator_2_io_out;
  wire [4:0] Accumulator_2_io_sel;
  wire  Accumulator_2_io_en;
  wire  Accumulator_2_io_reset;
  wire [3:0] _T_1275;
  wire [3:0] _T_1276;
  wire [3:0] _T_1277;
  wire [3:0] _T_1278;
  wire [3:0] _T_1279;
  wire [3:0] _T_1280;
  wire [3:0] _T_1281;
  wire [3:0] _T_1282;
  reg [5:0] _T_1285;
  reg [31:0] _GEN_772;
  reg [5:0] _T_1288;
  reg [31:0] _GEN_773;
  reg [5:0] _T_1291;
  reg [31:0] _GEN_774;
  reg [5:0] _T_1294;
  reg [31:0] _GEN_775;
  reg [5:0] _T_1297;
  reg [31:0] _GEN_776;
  reg [5:0] _T_1300;
  reg [31:0] _GEN_777;
  reg [5:0] _T_1303;
  reg [31:0] _GEN_778;
  reg [5:0] _T_1306;
  reg [31:0] _GEN_779;
  reg [5:0] _T_1309;
  reg [31:0] _GEN_780;
  reg [5:0] _T_1312;
  reg [31:0] _GEN_781;
  reg [5:0] _T_1315;
  reg [31:0] _GEN_782;
  reg [5:0] _T_1318;
  reg [31:0] _GEN_783;
  reg [5:0] _T_1321;
  reg [31:0] _GEN_784;
  reg [5:0] _T_1324;
  reg [31:0] _GEN_785;
  reg [5:0] _T_1327;
  reg [31:0] _GEN_786;
  reg [5:0] _T_1330;
  reg [31:0] _GEN_787;
  wire [5:0] _T_1333_0;
  wire [5:0] _T_1333_1;
  wire [5:0] _T_1333_2;
  wire [5:0] _T_1333_3;
  wire [5:0] _T_1333_4;
  wire [5:0] _T_1333_5;
  wire [5:0] _T_1333_6;
  wire [5:0] _T_1333_7;
  wire [5:0] _T_1333_8;
  wire [5:0] _T_1333_9;
  wire [5:0] _T_1333_10;
  wire [5:0] _T_1333_11;
  wire [5:0] _T_1333_12;
  wire [5:0] _T_1333_13;
  wire [5:0] _T_1333_14;
  wire [5:0] _T_1333_15;
  reg [5:0] _T_1355;
  reg [31:0] _GEN_788;
  reg [5:0] _T_1358;
  reg [31:0] _GEN_789;
  reg [5:0] _T_1361;
  reg [31:0] _GEN_790;
  reg [5:0] _T_1364;
  reg [31:0] _GEN_791;
  reg [5:0] _T_1367;
  reg [31:0] _GEN_792;
  reg [5:0] _T_1370;
  reg [31:0] _GEN_793;
  reg [5:0] _T_1373;
  reg [31:0] _GEN_794;
  reg [5:0] _T_1376;
  reg [31:0] _GEN_795;
  reg [5:0] _T_1379;
  reg [31:0] _GEN_796;
  reg [5:0] _T_1382;
  reg [31:0] _GEN_797;
  reg [5:0] _T_1385;
  reg [31:0] _GEN_798;
  reg [5:0] _T_1388;
  reg [31:0] _GEN_799;
  reg [5:0] _T_1391;
  reg [31:0] _GEN_800;
  reg [5:0] _T_1394;
  reg [31:0] _GEN_801;
  reg [5:0] _T_1397;
  reg [31:0] _GEN_802;
  reg [5:0] _T_1400;
  reg [31:0] _GEN_803;
  wire [5:0] _T_1403_0;
  wire [5:0] _T_1403_1;
  wire [5:0] _T_1403_2;
  wire [5:0] _T_1403_3;
  wire [5:0] _T_1403_4;
  wire [5:0] _T_1403_5;
  wire [5:0] _T_1403_6;
  wire [5:0] _T_1403_7;
  wire [5:0] _T_1403_8;
  wire [5:0] _T_1403_9;
  wire [5:0] _T_1403_10;
  wire [5:0] _T_1403_11;
  wire [5:0] _T_1403_12;
  wire [5:0] _T_1403_13;
  wire [5:0] _T_1403_14;
  wire [5:0] _T_1403_15;
  reg [5:0] _T_1425;
  reg [31:0] _GEN_804;
  reg [5:0] _T_1428;
  reg [31:0] _GEN_805;
  reg [5:0] _T_1431;
  reg [31:0] _GEN_806;
  reg [5:0] _T_1434;
  reg [31:0] _GEN_807;
  reg [5:0] _T_1437;
  reg [31:0] _GEN_808;
  reg [5:0] _T_1440;
  reg [31:0] _GEN_809;
  reg [5:0] _T_1443;
  reg [31:0] _GEN_810;
  reg [5:0] _T_1446;
  reg [31:0] _GEN_811;
  reg [5:0] _T_1449;
  reg [31:0] _GEN_812;
  reg [5:0] _T_1452;
  reg [31:0] _GEN_813;
  reg [5:0] _T_1455;
  reg [31:0] _GEN_814;
  reg [5:0] _T_1458;
  reg [31:0] _GEN_815;
  reg [5:0] _T_1461;
  reg [31:0] _GEN_816;
  reg [5:0] _T_1464;
  reg [31:0] _GEN_817;
  reg [5:0] _T_1467;
  reg [31:0] _GEN_818;
  reg [5:0] _T_1470;
  reg [31:0] _GEN_819;
  wire [5:0] _T_1473_0;
  wire [5:0] _T_1473_1;
  wire [5:0] _T_1473_2;
  wire [5:0] _T_1473_3;
  wire [5:0] _T_1473_4;
  wire [5:0] _T_1473_5;
  wire [5:0] _T_1473_6;
  wire [5:0] _T_1473_7;
  wire [5:0] _T_1473_8;
  wire [5:0] _T_1473_9;
  wire [5:0] _T_1473_10;
  wire [5:0] _T_1473_11;
  wire [5:0] _T_1473_12;
  wire [5:0] _T_1473_13;
  wire [5:0] _T_1473_14;
  wire [5:0] _T_1473_15;
  reg [5:0] _T_1495;
  reg [31:0] _GEN_820;
  reg [5:0] _T_1498;
  reg [31:0] _GEN_821;
  reg [5:0] _T_1501;
  reg [31:0] _GEN_822;
  reg [5:0] _T_1504;
  reg [31:0] _GEN_823;
  reg [5:0] _T_1507;
  reg [31:0] _GEN_824;
  reg [5:0] _T_1510;
  reg [31:0] _GEN_825;
  reg [5:0] _T_1513;
  reg [31:0] _GEN_826;
  reg [5:0] _T_1516;
  reg [31:0] _GEN_827;
  reg [5:0] _T_1519;
  reg [31:0] _GEN_828;
  reg [5:0] _T_1522;
  reg [31:0] _GEN_829;
  reg [5:0] _T_1525;
  reg [31:0] _GEN_830;
  reg [5:0] _T_1528;
  reg [31:0] _GEN_831;
  reg [5:0] _T_1531;
  reg [31:0] _GEN_832;
  reg [5:0] _T_1534;
  reg [31:0] _GEN_833;
  reg [5:0] _T_1537;
  reg [31:0] _GEN_834;
  reg [5:0] _T_1540;
  reg [31:0] _GEN_835;
  wire [5:0] _T_1543_0;
  wire [5:0] _T_1543_1;
  wire [5:0] _T_1543_2;
  wire [5:0] _T_1543_3;
  wire [5:0] _T_1543_4;
  wire [5:0] _T_1543_5;
  wire [5:0] _T_1543_6;
  wire [5:0] _T_1543_7;
  wire [5:0] _T_1543_8;
  wire [5:0] _T_1543_9;
  wire [5:0] _T_1543_10;
  wire [5:0] _T_1543_11;
  wire [5:0] _T_1543_12;
  wire [5:0] _T_1543_13;
  wire [5:0] _T_1543_14;
  wire [5:0] _T_1543_15;
  reg [5:0] _T_1565;
  reg [31:0] _GEN_836;
  reg [5:0] _T_1568;
  reg [31:0] _GEN_837;
  reg [5:0] _T_1571;
  reg [31:0] _GEN_838;
  reg [5:0] _T_1574;
  reg [31:0] _GEN_839;
  reg [5:0] _T_1577;
  reg [31:0] _GEN_840;
  reg [5:0] _T_1580;
  reg [31:0] _GEN_841;
  reg [5:0] _T_1583;
  reg [31:0] _GEN_842;
  reg [5:0] _T_1586;
  reg [31:0] _GEN_843;
  reg [5:0] _T_1589;
  reg [31:0] _GEN_844;
  reg [5:0] _T_1592;
  reg [31:0] _GEN_845;
  reg [5:0] _T_1595;
  reg [31:0] _GEN_846;
  reg [5:0] _T_1598;
  reg [31:0] _GEN_847;
  reg [5:0] _T_1601;
  reg [31:0] _GEN_848;
  reg [5:0] _T_1604;
  reg [31:0] _GEN_849;
  reg [5:0] _T_1607;
  reg [31:0] _GEN_850;
  reg [5:0] _T_1610;
  reg [31:0] _GEN_851;
  wire [5:0] _T_1613_0;
  wire [5:0] _T_1613_1;
  wire [5:0] _T_1613_2;
  wire [5:0] _T_1613_3;
  wire [5:0] _T_1613_4;
  wire [5:0] _T_1613_5;
  wire [5:0] _T_1613_6;
  wire [5:0] _T_1613_7;
  wire [5:0] _T_1613_8;
  wire [5:0] _T_1613_9;
  wire [5:0] _T_1613_10;
  wire [5:0] _T_1613_11;
  wire [5:0] _T_1613_12;
  wire [5:0] _T_1613_13;
  wire [5:0] _T_1613_14;
  wire [5:0] _T_1613_15;
  reg [5:0] _T_1635;
  reg [31:0] _GEN_852;
  reg [5:0] _T_1638;
  reg [31:0] _GEN_853;
  reg [5:0] _T_1641;
  reg [31:0] _GEN_854;
  reg [5:0] _T_1644;
  reg [31:0] _GEN_855;
  reg [5:0] _T_1647;
  reg [31:0] _GEN_856;
  reg [5:0] _T_1650;
  reg [31:0] _GEN_857;
  reg [5:0] _T_1653;
  reg [31:0] _GEN_858;
  reg [5:0] _T_1656;
  reg [31:0] _GEN_859;
  reg [5:0] _T_1659;
  reg [31:0] _GEN_860;
  reg [5:0] _T_1662;
  reg [31:0] _GEN_861;
  reg [5:0] _T_1665;
  reg [31:0] _GEN_862;
  reg [5:0] _T_1668;
  reg [31:0] _GEN_863;
  reg [5:0] _T_1671;
  reg [31:0] _GEN_864;
  reg [5:0] _T_1674;
  reg [31:0] _GEN_865;
  reg [5:0] _T_1677;
  reg [31:0] _GEN_866;
  reg [5:0] _T_1680;
  reg [31:0] _GEN_867;
  wire [5:0] _T_1683_0;
  wire [5:0] _T_1683_1;
  wire [5:0] _T_1683_2;
  wire [5:0] _T_1683_3;
  wire [5:0] _T_1683_4;
  wire [5:0] _T_1683_5;
  wire [5:0] _T_1683_6;
  wire [5:0] _T_1683_7;
  wire [5:0] _T_1683_8;
  wire [5:0] _T_1683_9;
  wire [5:0] _T_1683_10;
  wire [5:0] _T_1683_11;
  wire [5:0] _T_1683_12;
  wire [5:0] _T_1683_13;
  wire [5:0] _T_1683_14;
  wire [5:0] _T_1683_15;
  reg [5:0] _T_1705;
  reg [31:0] _GEN_868;
  reg [5:0] _T_1708;
  reg [31:0] _GEN_869;
  reg [5:0] _T_1711;
  reg [31:0] _GEN_870;
  reg [5:0] _T_1714;
  reg [31:0] _GEN_871;
  reg [5:0] _T_1717;
  reg [31:0] _GEN_872;
  reg [5:0] _T_1720;
  reg [31:0] _GEN_873;
  reg [5:0] _T_1723;
  reg [31:0] _GEN_874;
  reg [5:0] _T_1726;
  reg [31:0] _GEN_875;
  reg [5:0] _T_1729;
  reg [31:0] _GEN_876;
  reg [5:0] _T_1732;
  reg [31:0] _GEN_877;
  reg [5:0] _T_1735;
  reg [31:0] _GEN_878;
  reg [5:0] _T_1738;
  reg [31:0] _GEN_879;
  reg [5:0] _T_1741;
  reg [31:0] _GEN_880;
  reg [5:0] _T_1744;
  reg [31:0] _GEN_881;
  reg [5:0] _T_1747;
  reg [31:0] _GEN_882;
  reg [5:0] _T_1750;
  reg [31:0] _GEN_883;
  wire [5:0] _T_1753_0;
  wire [5:0] _T_1753_1;
  wire [5:0] _T_1753_2;
  wire [5:0] _T_1753_3;
  wire [5:0] _T_1753_4;
  wire [5:0] _T_1753_5;
  wire [5:0] _T_1753_6;
  wire [5:0] _T_1753_7;
  wire [5:0] _T_1753_8;
  wire [5:0] _T_1753_9;
  wire [5:0] _T_1753_10;
  wire [5:0] _T_1753_11;
  wire [5:0] _T_1753_12;
  wire [5:0] _T_1753_13;
  wire [5:0] _T_1753_14;
  wire [5:0] _T_1753_15;
  reg [5:0] _T_1775;
  reg [31:0] _GEN_884;
  reg [5:0] _T_1778;
  reg [31:0] _GEN_885;
  reg [5:0] _T_1781;
  reg [31:0] _GEN_886;
  reg [5:0] _T_1784;
  reg [31:0] _GEN_887;
  reg [5:0] _T_1787;
  reg [31:0] _GEN_888;
  reg [5:0] _T_1790;
  reg [31:0] _GEN_889;
  reg [5:0] _T_1793;
  reg [31:0] _GEN_890;
  reg [5:0] _T_1796;
  reg [31:0] _GEN_891;
  reg [5:0] _T_1799;
  reg [31:0] _GEN_892;
  reg [5:0] _T_1802;
  reg [31:0] _GEN_893;
  reg [5:0] _T_1805;
  reg [31:0] _GEN_894;
  reg [5:0] _T_1808;
  reg [31:0] _GEN_895;
  reg [5:0] _T_1811;
  reg [31:0] _GEN_896;
  reg [5:0] _T_1814;
  reg [31:0] _GEN_897;
  reg [5:0] _T_1817;
  reg [31:0] _GEN_898;
  reg [5:0] _T_1820;
  reg [31:0] _GEN_899;
  wire [5:0] _T_1823_0;
  wire [5:0] _T_1823_1;
  wire [5:0] _T_1823_2;
  wire [5:0] _T_1823_3;
  wire [5:0] _T_1823_4;
  wire [5:0] _T_1823_5;
  wire [5:0] _T_1823_6;
  wire [5:0] _T_1823_7;
  wire [5:0] _T_1823_8;
  wire [5:0] _T_1823_9;
  wire [5:0] _T_1823_10;
  wire [5:0] _T_1823_11;
  wire [5:0] _T_1823_12;
  wire [5:0] _T_1823_13;
  wire [5:0] _T_1823_14;
  wire [5:0] _T_1823_15;
  wire [5:0] _GEN_16;
  wire [5:0] _GEN_272;
  wire [5:0] _GEN_273;
  wire [5:0] _GEN_274;
  wire [5:0] _GEN_275;
  wire [5:0] _GEN_276;
  wire [5:0] _GEN_277;
  wire [5:0] _GEN_278;
  wire [5:0] _GEN_279;
  wire [5:0] _GEN_280;
  wire [5:0] _GEN_281;
  wire [5:0] _GEN_282;
  wire [5:0] _GEN_283;
  wire [5:0] _GEN_284;
  wire [5:0] _GEN_285;
  wire [5:0] _GEN_286;
  wire [5:0] _GEN_17;
  wire [5:0] _GEN_287;
  wire [5:0] _GEN_288;
  wire [5:0] _GEN_289;
  wire [5:0] _GEN_290;
  wire [5:0] _GEN_291;
  wire [5:0] _GEN_292;
  wire [5:0] _GEN_293;
  wire [5:0] _GEN_294;
  wire [5:0] _GEN_295;
  wire [5:0] _GEN_296;
  wire [5:0] _GEN_297;
  wire [5:0] _GEN_298;
  wire [5:0] _GEN_299;
  wire [5:0] _GEN_300;
  wire [5:0] _GEN_301;
  wire [6:0] _T_1843;
  wire [5:0] _T_1844;
  wire [5:0] _T_1845;
  wire [5:0] _GEN_18;
  wire [5:0] _GEN_302;
  wire [5:0] _GEN_303;
  wire [5:0] _GEN_304;
  wire [5:0] _GEN_305;
  wire [5:0] _GEN_306;
  wire [5:0] _GEN_307;
  wire [5:0] _GEN_308;
  wire [5:0] _GEN_309;
  wire [5:0] _GEN_310;
  wire [5:0] _GEN_311;
  wire [5:0] _GEN_312;
  wire [5:0] _GEN_313;
  wire [5:0] _GEN_314;
  wire [5:0] _GEN_315;
  wire [5:0] _GEN_316;
  wire [5:0] _GEN_19;
  wire [5:0] _GEN_317;
  wire [5:0] _GEN_318;
  wire [5:0] _GEN_319;
  wire [5:0] _GEN_320;
  wire [5:0] _GEN_321;
  wire [5:0] _GEN_322;
  wire [5:0] _GEN_323;
  wire [5:0] _GEN_324;
  wire [5:0] _GEN_325;
  wire [5:0] _GEN_326;
  wire [5:0] _GEN_327;
  wire [5:0] _GEN_328;
  wire [5:0] _GEN_329;
  wire [5:0] _GEN_330;
  wire [5:0] _GEN_331;
  wire [6:0] _T_1846;
  wire [5:0] _T_1847;
  wire [5:0] _T_1848;
  wire [5:0] _GEN_20;
  wire [5:0] _GEN_332;
  wire [5:0] _GEN_333;
  wire [5:0] _GEN_334;
  wire [5:0] _GEN_335;
  wire [5:0] _GEN_336;
  wire [5:0] _GEN_337;
  wire [5:0] _GEN_338;
  wire [5:0] _GEN_339;
  wire [5:0] _GEN_340;
  wire [5:0] _GEN_341;
  wire [5:0] _GEN_342;
  wire [5:0] _GEN_343;
  wire [5:0] _GEN_344;
  wire [5:0] _GEN_345;
  wire [5:0] _GEN_346;
  wire [5:0] _GEN_21;
  wire [5:0] _GEN_347;
  wire [5:0] _GEN_348;
  wire [5:0] _GEN_349;
  wire [5:0] _GEN_350;
  wire [5:0] _GEN_351;
  wire [5:0] _GEN_352;
  wire [5:0] _GEN_353;
  wire [5:0] _GEN_354;
  wire [5:0] _GEN_355;
  wire [5:0] _GEN_356;
  wire [5:0] _GEN_357;
  wire [5:0] _GEN_358;
  wire [5:0] _GEN_359;
  wire [5:0] _GEN_360;
  wire [5:0] _GEN_361;
  wire [6:0] _T_1849;
  wire [5:0] _T_1850;
  wire [5:0] _T_1851;
  wire [5:0] _GEN_22;
  wire [5:0] _GEN_362;
  wire [5:0] _GEN_363;
  wire [5:0] _GEN_364;
  wire [5:0] _GEN_365;
  wire [5:0] _GEN_366;
  wire [5:0] _GEN_367;
  wire [5:0] _GEN_368;
  wire [5:0] _GEN_369;
  wire [5:0] _GEN_370;
  wire [5:0] _GEN_371;
  wire [5:0] _GEN_372;
  wire [5:0] _GEN_373;
  wire [5:0] _GEN_374;
  wire [5:0] _GEN_375;
  wire [5:0] _GEN_376;
  wire [5:0] _GEN_23;
  wire [5:0] _GEN_377;
  wire [5:0] _GEN_378;
  wire [5:0] _GEN_379;
  wire [5:0] _GEN_380;
  wire [5:0] _GEN_381;
  wire [5:0] _GEN_382;
  wire [5:0] _GEN_383;
  wire [5:0] _GEN_384;
  wire [5:0] _GEN_385;
  wire [5:0] _GEN_386;
  wire [5:0] _GEN_387;
  wire [5:0] _GEN_388;
  wire [5:0] _GEN_389;
  wire [5:0] _GEN_390;
  wire [5:0] _GEN_391;
  wire [6:0] _T_1852;
  wire [5:0] _T_1853;
  wire [5:0] _T_1854;
  wire [6:0] _T_1855;
  wire [5:0] _T_1856;
  wire [5:0] _T_1857;
  wire [6:0] _T_1858;
  wire [5:0] _T_1859;
  wire [5:0] _T_1860;
  wire [6:0] _T_1861;
  wire [5:0] _T_1862;
  wire [5:0] _T_1863;
  wire [15:0] MulAdd_2_io_a;
  wire [15:0] MulAdd_2_io_b;
  wire [31:0] MulAdd_2_io_m;
  wire [15:0] MulAdd_2_io_c;
  wire [31:0] MulAdd_2_io_r;
  wire [31:0] _T_1865;
  wire [31:0] _T_1866;
  wire [15:0] _T_1867;
  wire [15:0] _T_1868;
  wire [15:0] _T_1869;
  wire [15:0] _T_1870;
  wire  signs_2;
  wire  Accumulator_3_clock;
  wire [31:0] Accumulator_3_io_in;
  wire [31:0] Accumulator_3_io_out;
  wire [4:0] Accumulator_3_io_sel;
  wire  Accumulator_3_io_en;
  wire  Accumulator_3_io_reset;
  wire [3:0] _T_1871;
  wire [3:0] _T_1872;
  wire [3:0] _T_1873;
  wire [3:0] _T_1874;
  wire [3:0] _T_1875;
  wire [3:0] _T_1876;
  wire [3:0] _T_1877;
  wire [3:0] _T_1878;
  reg [5:0] _T_1881;
  reg [31:0] _GEN_900;
  reg [5:0] _T_1884;
  reg [31:0] _GEN_901;
  reg [5:0] _T_1887;
  reg [31:0] _GEN_902;
  reg [5:0] _T_1890;
  reg [31:0] _GEN_903;
  reg [5:0] _T_1893;
  reg [31:0] _GEN_904;
  reg [5:0] _T_1896;
  reg [31:0] _GEN_905;
  reg [5:0] _T_1899;
  reg [31:0] _GEN_906;
  reg [5:0] _T_1902;
  reg [31:0] _GEN_907;
  reg [5:0] _T_1905;
  reg [31:0] _GEN_908;
  reg [5:0] _T_1908;
  reg [31:0] _GEN_909;
  reg [5:0] _T_1911;
  reg [31:0] _GEN_910;
  reg [5:0] _T_1914;
  reg [31:0] _GEN_911;
  reg [5:0] _T_1917;
  reg [31:0] _GEN_912;
  reg [5:0] _T_1920;
  reg [31:0] _GEN_913;
  reg [5:0] _T_1923;
  reg [31:0] _GEN_914;
  reg [5:0] _T_1926;
  reg [31:0] _GEN_915;
  wire [5:0] _T_1929_0;
  wire [5:0] _T_1929_1;
  wire [5:0] _T_1929_2;
  wire [5:0] _T_1929_3;
  wire [5:0] _T_1929_4;
  wire [5:0] _T_1929_5;
  wire [5:0] _T_1929_6;
  wire [5:0] _T_1929_7;
  wire [5:0] _T_1929_8;
  wire [5:0] _T_1929_9;
  wire [5:0] _T_1929_10;
  wire [5:0] _T_1929_11;
  wire [5:0] _T_1929_12;
  wire [5:0] _T_1929_13;
  wire [5:0] _T_1929_14;
  wire [5:0] _T_1929_15;
  reg [5:0] _T_1951;
  reg [31:0] _GEN_916;
  reg [5:0] _T_1954;
  reg [31:0] _GEN_917;
  reg [5:0] _T_1957;
  reg [31:0] _GEN_918;
  reg [5:0] _T_1960;
  reg [31:0] _GEN_919;
  reg [5:0] _T_1963;
  reg [31:0] _GEN_920;
  reg [5:0] _T_1966;
  reg [31:0] _GEN_921;
  reg [5:0] _T_1969;
  reg [31:0] _GEN_922;
  reg [5:0] _T_1972;
  reg [31:0] _GEN_923;
  reg [5:0] _T_1975;
  reg [31:0] _GEN_924;
  reg [5:0] _T_1978;
  reg [31:0] _GEN_925;
  reg [5:0] _T_1981;
  reg [31:0] _GEN_926;
  reg [5:0] _T_1984;
  reg [31:0] _GEN_927;
  reg [5:0] _T_1987;
  reg [31:0] _GEN_928;
  reg [5:0] _T_1990;
  reg [31:0] _GEN_929;
  reg [5:0] _T_1993;
  reg [31:0] _GEN_930;
  reg [5:0] _T_1996;
  reg [31:0] _GEN_931;
  wire [5:0] _T_1999_0;
  wire [5:0] _T_1999_1;
  wire [5:0] _T_1999_2;
  wire [5:0] _T_1999_3;
  wire [5:0] _T_1999_4;
  wire [5:0] _T_1999_5;
  wire [5:0] _T_1999_6;
  wire [5:0] _T_1999_7;
  wire [5:0] _T_1999_8;
  wire [5:0] _T_1999_9;
  wire [5:0] _T_1999_10;
  wire [5:0] _T_1999_11;
  wire [5:0] _T_1999_12;
  wire [5:0] _T_1999_13;
  wire [5:0] _T_1999_14;
  wire [5:0] _T_1999_15;
  reg [5:0] _T_2021;
  reg [31:0] _GEN_932;
  reg [5:0] _T_2024;
  reg [31:0] _GEN_933;
  reg [5:0] _T_2027;
  reg [31:0] _GEN_934;
  reg [5:0] _T_2030;
  reg [31:0] _GEN_935;
  reg [5:0] _T_2033;
  reg [31:0] _GEN_936;
  reg [5:0] _T_2036;
  reg [31:0] _GEN_937;
  reg [5:0] _T_2039;
  reg [31:0] _GEN_938;
  reg [5:0] _T_2042;
  reg [31:0] _GEN_939;
  reg [5:0] _T_2045;
  reg [31:0] _GEN_940;
  reg [5:0] _T_2048;
  reg [31:0] _GEN_941;
  reg [5:0] _T_2051;
  reg [31:0] _GEN_942;
  reg [5:0] _T_2054;
  reg [31:0] _GEN_943;
  reg [5:0] _T_2057;
  reg [31:0] _GEN_944;
  reg [5:0] _T_2060;
  reg [31:0] _GEN_945;
  reg [5:0] _T_2063;
  reg [31:0] _GEN_946;
  reg [5:0] _T_2066;
  reg [31:0] _GEN_947;
  wire [5:0] _T_2069_0;
  wire [5:0] _T_2069_1;
  wire [5:0] _T_2069_2;
  wire [5:0] _T_2069_3;
  wire [5:0] _T_2069_4;
  wire [5:0] _T_2069_5;
  wire [5:0] _T_2069_6;
  wire [5:0] _T_2069_7;
  wire [5:0] _T_2069_8;
  wire [5:0] _T_2069_9;
  wire [5:0] _T_2069_10;
  wire [5:0] _T_2069_11;
  wire [5:0] _T_2069_12;
  wire [5:0] _T_2069_13;
  wire [5:0] _T_2069_14;
  wire [5:0] _T_2069_15;
  reg [5:0] _T_2091;
  reg [31:0] _GEN_948;
  reg [5:0] _T_2094;
  reg [31:0] _GEN_949;
  reg [5:0] _T_2097;
  reg [31:0] _GEN_950;
  reg [5:0] _T_2100;
  reg [31:0] _GEN_951;
  reg [5:0] _T_2103;
  reg [31:0] _GEN_952;
  reg [5:0] _T_2106;
  reg [31:0] _GEN_953;
  reg [5:0] _T_2109;
  reg [31:0] _GEN_954;
  reg [5:0] _T_2112;
  reg [31:0] _GEN_955;
  reg [5:0] _T_2115;
  reg [31:0] _GEN_956;
  reg [5:0] _T_2118;
  reg [31:0] _GEN_957;
  reg [5:0] _T_2121;
  reg [31:0] _GEN_958;
  reg [5:0] _T_2124;
  reg [31:0] _GEN_959;
  reg [5:0] _T_2127;
  reg [31:0] _GEN_960;
  reg [5:0] _T_2130;
  reg [31:0] _GEN_961;
  reg [5:0] _T_2133;
  reg [31:0] _GEN_962;
  reg [5:0] _T_2136;
  reg [31:0] _GEN_963;
  wire [5:0] _T_2139_0;
  wire [5:0] _T_2139_1;
  wire [5:0] _T_2139_2;
  wire [5:0] _T_2139_3;
  wire [5:0] _T_2139_4;
  wire [5:0] _T_2139_5;
  wire [5:0] _T_2139_6;
  wire [5:0] _T_2139_7;
  wire [5:0] _T_2139_8;
  wire [5:0] _T_2139_9;
  wire [5:0] _T_2139_10;
  wire [5:0] _T_2139_11;
  wire [5:0] _T_2139_12;
  wire [5:0] _T_2139_13;
  wire [5:0] _T_2139_14;
  wire [5:0] _T_2139_15;
  reg [5:0] _T_2161;
  reg [31:0] _GEN_964;
  reg [5:0] _T_2164;
  reg [31:0] _GEN_965;
  reg [5:0] _T_2167;
  reg [31:0] _GEN_966;
  reg [5:0] _T_2170;
  reg [31:0] _GEN_967;
  reg [5:0] _T_2173;
  reg [31:0] _GEN_968;
  reg [5:0] _T_2176;
  reg [31:0] _GEN_969;
  reg [5:0] _T_2179;
  reg [31:0] _GEN_970;
  reg [5:0] _T_2182;
  reg [31:0] _GEN_971;
  reg [5:0] _T_2185;
  reg [31:0] _GEN_972;
  reg [5:0] _T_2188;
  reg [31:0] _GEN_973;
  reg [5:0] _T_2191;
  reg [31:0] _GEN_974;
  reg [5:0] _T_2194;
  reg [31:0] _GEN_975;
  reg [5:0] _T_2197;
  reg [31:0] _GEN_976;
  reg [5:0] _T_2200;
  reg [31:0] _GEN_977;
  reg [5:0] _T_2203;
  reg [31:0] _GEN_978;
  reg [5:0] _T_2206;
  reg [31:0] _GEN_979;
  wire [5:0] _T_2209_0;
  wire [5:0] _T_2209_1;
  wire [5:0] _T_2209_2;
  wire [5:0] _T_2209_3;
  wire [5:0] _T_2209_4;
  wire [5:0] _T_2209_5;
  wire [5:0] _T_2209_6;
  wire [5:0] _T_2209_7;
  wire [5:0] _T_2209_8;
  wire [5:0] _T_2209_9;
  wire [5:0] _T_2209_10;
  wire [5:0] _T_2209_11;
  wire [5:0] _T_2209_12;
  wire [5:0] _T_2209_13;
  wire [5:0] _T_2209_14;
  wire [5:0] _T_2209_15;
  reg [5:0] _T_2231;
  reg [31:0] _GEN_980;
  reg [5:0] _T_2234;
  reg [31:0] _GEN_981;
  reg [5:0] _T_2237;
  reg [31:0] _GEN_982;
  reg [5:0] _T_2240;
  reg [31:0] _GEN_983;
  reg [5:0] _T_2243;
  reg [31:0] _GEN_984;
  reg [5:0] _T_2246;
  reg [31:0] _GEN_985;
  reg [5:0] _T_2249;
  reg [31:0] _GEN_986;
  reg [5:0] _T_2252;
  reg [31:0] _GEN_987;
  reg [5:0] _T_2255;
  reg [31:0] _GEN_988;
  reg [5:0] _T_2258;
  reg [31:0] _GEN_989;
  reg [5:0] _T_2261;
  reg [31:0] _GEN_990;
  reg [5:0] _T_2264;
  reg [31:0] _GEN_991;
  reg [5:0] _T_2267;
  reg [31:0] _GEN_992;
  reg [5:0] _T_2270;
  reg [31:0] _GEN_993;
  reg [5:0] _T_2273;
  reg [31:0] _GEN_994;
  reg [5:0] _T_2276;
  reg [31:0] _GEN_995;
  wire [5:0] _T_2279_0;
  wire [5:0] _T_2279_1;
  wire [5:0] _T_2279_2;
  wire [5:0] _T_2279_3;
  wire [5:0] _T_2279_4;
  wire [5:0] _T_2279_5;
  wire [5:0] _T_2279_6;
  wire [5:0] _T_2279_7;
  wire [5:0] _T_2279_8;
  wire [5:0] _T_2279_9;
  wire [5:0] _T_2279_10;
  wire [5:0] _T_2279_11;
  wire [5:0] _T_2279_12;
  wire [5:0] _T_2279_13;
  wire [5:0] _T_2279_14;
  wire [5:0] _T_2279_15;
  reg [5:0] _T_2301;
  reg [31:0] _GEN_996;
  reg [5:0] _T_2304;
  reg [31:0] _GEN_997;
  reg [5:0] _T_2307;
  reg [31:0] _GEN_998;
  reg [5:0] _T_2310;
  reg [31:0] _GEN_999;
  reg [5:0] _T_2313;
  reg [31:0] _GEN_1000;
  reg [5:0] _T_2316;
  reg [31:0] _GEN_1001;
  reg [5:0] _T_2319;
  reg [31:0] _GEN_1002;
  reg [5:0] _T_2322;
  reg [31:0] _GEN_1003;
  reg [5:0] _T_2325;
  reg [31:0] _GEN_1004;
  reg [5:0] _T_2328;
  reg [31:0] _GEN_1005;
  reg [5:0] _T_2331;
  reg [31:0] _GEN_1006;
  reg [5:0] _T_2334;
  reg [31:0] _GEN_1007;
  reg [5:0] _T_2337;
  reg [31:0] _GEN_1008;
  reg [5:0] _T_2340;
  reg [31:0] _GEN_1009;
  reg [5:0] _T_2343;
  reg [31:0] _GEN_1010;
  reg [5:0] _T_2346;
  reg [31:0] _GEN_1011;
  wire [5:0] _T_2349_0;
  wire [5:0] _T_2349_1;
  wire [5:0] _T_2349_2;
  wire [5:0] _T_2349_3;
  wire [5:0] _T_2349_4;
  wire [5:0] _T_2349_5;
  wire [5:0] _T_2349_6;
  wire [5:0] _T_2349_7;
  wire [5:0] _T_2349_8;
  wire [5:0] _T_2349_9;
  wire [5:0] _T_2349_10;
  wire [5:0] _T_2349_11;
  wire [5:0] _T_2349_12;
  wire [5:0] _T_2349_13;
  wire [5:0] _T_2349_14;
  wire [5:0] _T_2349_15;
  reg [5:0] _T_2371;
  reg [31:0] _GEN_1012;
  reg [5:0] _T_2374;
  reg [31:0] _GEN_1013;
  reg [5:0] _T_2377;
  reg [31:0] _GEN_1014;
  reg [5:0] _T_2380;
  reg [31:0] _GEN_1015;
  reg [5:0] _T_2383;
  reg [31:0] _GEN_1016;
  reg [5:0] _T_2386;
  reg [31:0] _GEN_1017;
  reg [5:0] _T_2389;
  reg [31:0] _GEN_1018;
  reg [5:0] _T_2392;
  reg [31:0] _GEN_1019;
  reg [5:0] _T_2395;
  reg [31:0] _GEN_1020;
  reg [5:0] _T_2398;
  reg [31:0] _GEN_1021;
  reg [5:0] _T_2401;
  reg [31:0] _GEN_1022;
  reg [5:0] _T_2404;
  reg [31:0] _GEN_1023;
  reg [5:0] _T_2407;
  reg [31:0] _GEN_1024;
  reg [5:0] _T_2410;
  reg [31:0] _GEN_1025;
  reg [5:0] _T_2413;
  reg [31:0] _GEN_1026;
  reg [5:0] _T_2416;
  reg [31:0] _GEN_1027;
  wire [5:0] _T_2419_0;
  wire [5:0] _T_2419_1;
  wire [5:0] _T_2419_2;
  wire [5:0] _T_2419_3;
  wire [5:0] _T_2419_4;
  wire [5:0] _T_2419_5;
  wire [5:0] _T_2419_6;
  wire [5:0] _T_2419_7;
  wire [5:0] _T_2419_8;
  wire [5:0] _T_2419_9;
  wire [5:0] _T_2419_10;
  wire [5:0] _T_2419_11;
  wire [5:0] _T_2419_12;
  wire [5:0] _T_2419_13;
  wire [5:0] _T_2419_14;
  wire [5:0] _T_2419_15;
  wire [5:0] _GEN_24;
  wire [5:0] _GEN_392;
  wire [5:0] _GEN_393;
  wire [5:0] _GEN_394;
  wire [5:0] _GEN_395;
  wire [5:0] _GEN_396;
  wire [5:0] _GEN_397;
  wire [5:0] _GEN_398;
  wire [5:0] _GEN_399;
  wire [5:0] _GEN_400;
  wire [5:0] _GEN_401;
  wire [5:0] _GEN_402;
  wire [5:0] _GEN_403;
  wire [5:0] _GEN_404;
  wire [5:0] _GEN_405;
  wire [5:0] _GEN_406;
  wire [5:0] _GEN_25;
  wire [5:0] _GEN_407;
  wire [5:0] _GEN_408;
  wire [5:0] _GEN_409;
  wire [5:0] _GEN_410;
  wire [5:0] _GEN_411;
  wire [5:0] _GEN_412;
  wire [5:0] _GEN_413;
  wire [5:0] _GEN_414;
  wire [5:0] _GEN_415;
  wire [5:0] _GEN_416;
  wire [5:0] _GEN_417;
  wire [5:0] _GEN_418;
  wire [5:0] _GEN_419;
  wire [5:0] _GEN_420;
  wire [5:0] _GEN_421;
  wire [6:0] _T_2439;
  wire [5:0] _T_2440;
  wire [5:0] _T_2441;
  wire [5:0] _GEN_26;
  wire [5:0] _GEN_422;
  wire [5:0] _GEN_423;
  wire [5:0] _GEN_424;
  wire [5:0] _GEN_425;
  wire [5:0] _GEN_426;
  wire [5:0] _GEN_427;
  wire [5:0] _GEN_428;
  wire [5:0] _GEN_429;
  wire [5:0] _GEN_430;
  wire [5:0] _GEN_431;
  wire [5:0] _GEN_432;
  wire [5:0] _GEN_433;
  wire [5:0] _GEN_434;
  wire [5:0] _GEN_435;
  wire [5:0] _GEN_436;
  wire [5:0] _GEN_27;
  wire [5:0] _GEN_437;
  wire [5:0] _GEN_438;
  wire [5:0] _GEN_439;
  wire [5:0] _GEN_440;
  wire [5:0] _GEN_441;
  wire [5:0] _GEN_442;
  wire [5:0] _GEN_443;
  wire [5:0] _GEN_444;
  wire [5:0] _GEN_445;
  wire [5:0] _GEN_446;
  wire [5:0] _GEN_447;
  wire [5:0] _GEN_448;
  wire [5:0] _GEN_449;
  wire [5:0] _GEN_450;
  wire [5:0] _GEN_451;
  wire [6:0] _T_2442;
  wire [5:0] _T_2443;
  wire [5:0] _T_2444;
  wire [5:0] _GEN_28;
  wire [5:0] _GEN_452;
  wire [5:0] _GEN_453;
  wire [5:0] _GEN_454;
  wire [5:0] _GEN_455;
  wire [5:0] _GEN_456;
  wire [5:0] _GEN_457;
  wire [5:0] _GEN_458;
  wire [5:0] _GEN_459;
  wire [5:0] _GEN_460;
  wire [5:0] _GEN_461;
  wire [5:0] _GEN_462;
  wire [5:0] _GEN_463;
  wire [5:0] _GEN_464;
  wire [5:0] _GEN_465;
  wire [5:0] _GEN_466;
  wire [5:0] _GEN_29;
  wire [5:0] _GEN_467;
  wire [5:0] _GEN_468;
  wire [5:0] _GEN_469;
  wire [5:0] _GEN_470;
  wire [5:0] _GEN_471;
  wire [5:0] _GEN_472;
  wire [5:0] _GEN_473;
  wire [5:0] _GEN_474;
  wire [5:0] _GEN_475;
  wire [5:0] _GEN_476;
  wire [5:0] _GEN_477;
  wire [5:0] _GEN_478;
  wire [5:0] _GEN_479;
  wire [5:0] _GEN_480;
  wire [5:0] _GEN_481;
  wire [6:0] _T_2445;
  wire [5:0] _T_2446;
  wire [5:0] _T_2447;
  wire [5:0] _GEN_30;
  wire [5:0] _GEN_482;
  wire [5:0] _GEN_483;
  wire [5:0] _GEN_484;
  wire [5:0] _GEN_485;
  wire [5:0] _GEN_486;
  wire [5:0] _GEN_487;
  wire [5:0] _GEN_488;
  wire [5:0] _GEN_489;
  wire [5:0] _GEN_490;
  wire [5:0] _GEN_491;
  wire [5:0] _GEN_492;
  wire [5:0] _GEN_493;
  wire [5:0] _GEN_494;
  wire [5:0] _GEN_495;
  wire [5:0] _GEN_496;
  wire [5:0] _GEN_31;
  wire [5:0] _GEN_497;
  wire [5:0] _GEN_498;
  wire [5:0] _GEN_499;
  wire [5:0] _GEN_500;
  wire [5:0] _GEN_501;
  wire [5:0] _GEN_502;
  wire [5:0] _GEN_503;
  wire [5:0] _GEN_504;
  wire [5:0] _GEN_505;
  wire [5:0] _GEN_506;
  wire [5:0] _GEN_507;
  wire [5:0] _GEN_508;
  wire [5:0] _GEN_509;
  wire [5:0] _GEN_510;
  wire [5:0] _GEN_511;
  wire [6:0] _T_2448;
  wire [5:0] _T_2449;
  wire [5:0] _T_2450;
  wire [6:0] _T_2451;
  wire [5:0] _T_2452;
  wire [5:0] _T_2453;
  wire [6:0] _T_2454;
  wire [5:0] _T_2455;
  wire [5:0] _T_2456;
  wire [6:0] _T_2457;
  wire [5:0] _T_2458;
  wire [5:0] _T_2459;
  wire [15:0] MulAdd_3_io_a;
  wire [15:0] MulAdd_3_io_b;
  wire [31:0] MulAdd_3_io_m;
  wire [15:0] MulAdd_3_io_c;
  wire [31:0] MulAdd_3_io_r;
  wire [31:0] _T_2461;
  wire [31:0] _T_2462;
  wire [15:0] _T_2463;
  wire [15:0] _T_2464;
  wire [15:0] _T_2465;
  wire [15:0] _T_2466;
  wire  signs_3;
  wire [1:0] _T_2467;
  wire [1:0] _T_2468;
  wire [3:0] _T_2469;
  wire [15:0] _GEN_512;
  wire [15:0] _GEN_513;
  wire [15:0] _GEN_514;
  wire [15:0] _GEN_515;
  AggregateMem mem (
    .clock(mem_clock),
    .io_addr(mem_io_addr),
    .io_in(mem_io_in),
    .io_out(mem_io_out),
    .io_wen(mem_io_wen),
    .io_ren(mem_io_ren)
  );
  BinaryBuffer binaryBuffer (
    .clock(binaryBuffer_clock),
    .reset(binaryBuffer_reset),
    .io_in(binaryBuffer_io_in),
    .io_push(binaryBuffer_io_push),
    .io_out(binaryBuffer_io_out),
    .io_pop(binaryBuffer_io_pop)
  );
  XNOR xnor$ (
    .io_in1(xnor$_io_in1),
    .io_in2_0(xnor$_io_in2_0),
    .io_in2_1(xnor$_io_in2_1),
    .io_in2_2(xnor$_io_in2_2),
    .io_in2_3(xnor$_io_in2_3),
    .io_out_0(xnor$_io_out_0),
    .io_out_1(xnor$_io_out_1),
    .io_out_2(xnor$_io_out_2),
    .io_out_3(xnor$_io_out_3)
  );
  MeanBuffer meanBuffer (
    .clock(meanBuffer_clock),
    .reset(meanBuffer_reset),
    .io_in_0(meanBuffer_io_in_0),
    .io_in_1(meanBuffer_io_in_1),
    .io_in_2(meanBuffer_io_in_2),
    .io_in_3(meanBuffer_io_in_3),
    .io_cntInverse65536(meanBuffer_io_cntInverse65536),
    .io_reset(meanBuffer_io_reset),
    .io_out(meanBuffer_io_out)
  );
  DelayedOutput mean (
    .clock(mean_clock),
    .reset(mean_reset),
    .io_input(mean_io_input),
    .io_update(mean_io_update),
    .io_output(mean_io_output)
  );
  MaxBuffer maxModule (
    .clock(maxModule_clock),
    .io_reset(maxModule_io_reset),
    .io_en(maxModule_io_en),
    .io_in_0(maxModule_io_in_0),
    .io_in_1(maxModule_io_in_1),
    .io_in_2(maxModule_io_in_2),
    .io_in_3(maxModule_io_in_3),
    .io_offset(maxModule_io_offset),
    .io_out(maxModule_io_out)
  );
  Accumulator Accumulator (
    .clock(Accumulator_clock),
    .io_in(Accumulator_io_in),
    .io_out(Accumulator_io_out),
    .io_sel(Accumulator_io_sel),
    .io_en(Accumulator_io_en),
    .io_reset(Accumulator_io_reset)
  );
  MulAdd MulAdd (
    .io_a(MulAdd_io_a),
    .io_b(MulAdd_io_b),
    .io_m(MulAdd_io_m),
    .io_c(MulAdd_io_c),
    .io_r(MulAdd_io_r)
  );
  Accumulator Accumulator_1 (
    .clock(Accumulator_1_clock),
    .io_in(Accumulator_1_io_in),
    .io_out(Accumulator_1_io_out),
    .io_sel(Accumulator_1_io_sel),
    .io_en(Accumulator_1_io_en),
    .io_reset(Accumulator_1_io_reset)
  );
  MulAdd MulAdd_1 (
    .io_a(MulAdd_1_io_a),
    .io_b(MulAdd_1_io_b),
    .io_m(MulAdd_1_io_m),
    .io_c(MulAdd_1_io_c),
    .io_r(MulAdd_1_io_r)
  );
  Accumulator Accumulator_2 (
    .clock(Accumulator_2_clock),
    .io_in(Accumulator_2_io_in),
    .io_out(Accumulator_2_io_out),
    .io_sel(Accumulator_2_io_sel),
    .io_en(Accumulator_2_io_en),
    .io_reset(Accumulator_2_io_reset)
  );
  MulAdd MulAdd_2 (
    .io_a(MulAdd_2_io_a),
    .io_b(MulAdd_2_io_b),
    .io_m(MulAdd_2_io_m),
    .io_c(MulAdd_2_io_c),
    .io_r(MulAdd_2_io_r)
  );
  Accumulator Accumulator_3 (
    .clock(Accumulator_3_clock),
    .io_in(Accumulator_3_io_in),
    .io_out(Accumulator_3_io_out),
    .io_sel(Accumulator_3_io_sel),
    .io_en(Accumulator_3_io_en),
    .io_reset(Accumulator_3_io_reset)
  );
  MulAdd MulAdd_3 (
    .io_a(MulAdd_3_io_a),
    .io_b(MulAdd_3_io_b),
    .io_m(MulAdd_3_io_m),
    .io_c(MulAdd_3_io_c),
    .io_r(MulAdd_3_io_r)
  );
  assign io_memOut = mem_io_out;
  assign io_result = maxModule_io_out;
  assign mem_clock = clock;
  assign mem_io_addr = io_memAddr;
  assign mem_io_in = io_memIn;
  assign mem_io_wen = io_memWen;
  assign mem_io_ren = io_memRen;
  assign inputWire = _T_2469;
  assign binaryBuffer_clock = clock;
  assign binaryBuffer_reset = reset;
  assign binaryBuffer_io_in = _T_24;
  assign binaryBuffer_io_push = io_inputBufferPush;
  assign binaryBuffer_io_pop = io_inputBufferPop;
  assign _T_24 = io_inputSel ? io_input : inputWire;
  assign xnor$_io_in1 = binaryBuffer_io_out;
  assign xnor$_io_in2_0 = _T_66_0;
  assign xnor$_io_in2_1 = _T_66_1;
  assign xnor$_io_in2_2 = _T_66_2;
  assign xnor$_io_in2_3 = _T_66_3;
  assign _T_35_0 = _T_49;
  assign _T_35_1 = _T_50;
  assign _T_35_2 = _T_51;
  assign _T_35_3 = _T_52;
  assign _T_48 = mem_io_out;
  assign _T_49 = _T_48[31:0];
  assign _T_50 = _T_48[63:32];
  assign _T_51 = _T_48[95:64];
  assign _T_52 = _T_48[127:96];
  assign _T_59_0 = 32'h0;
  assign _T_59_1 = 32'h0;
  assign _T_59_2 = 32'h0;
  assign _T_59_3 = 32'h0;
  assign _T_66_0 = io_memSel ? _T_35_0 : _T_59_0;
  assign _T_66_1 = io_memSel ? _T_35_1 : _T_59_1;
  assign _T_66_2 = io_memSel ? _T_35_2 : _T_59_2;
  assign _T_66_3 = io_memSel ? _T_35_3 : _T_59_3;
  assign meanBuffer_clock = clock;
  assign meanBuffer_reset = reset;
  assign meanBuffer_io_in_0 = MulAdd_io_r;
  assign meanBuffer_io_in_1 = MulAdd_1_io_r;
  assign meanBuffer_io_in_2 = MulAdd_2_io_r;
  assign meanBuffer_io_in_3 = MulAdd_3_io_r;
  assign meanBuffer_io_cntInverse65536 = io_featureNumInverse65536;
  assign meanBuffer_io_reset = io_meanReset;
  assign mean_clock = clock;
  assign mean_reset = reset;
  assign mean_io_input = meanBuffer_io_out;
  assign mean_io_update = io_meanUpdate;
  assign maxModule_clock = clock;
  assign maxModule_io_reset = io_maxClear;
  assign maxModule_io_en = io_maxEn;
  assign maxModule_io_in_0 = MulAdd_io_r;
  assign maxModule_io_in_1 = MulAdd_1_io_r;
  assign maxModule_io_in_2 = MulAdd_2_io_r;
  assign maxModule_io_in_3 = MulAdd_3_io_r;
  assign maxModule_io_offset = io_maxOffset;
  assign Accumulator_clock = clock;
  assign Accumulator_io_in = {{26{_T_671[5]}},_T_671};
  assign Accumulator_io_sel = io_accSel;
  assign Accumulator_io_en = io_accEn;
  assign Accumulator_io_reset = io_accReset;
  assign _T_83 = xnor$_io_out_0[3:0];
  assign _T_84 = xnor$_io_out_0[7:4];
  assign _T_85 = xnor$_io_out_0[11:8];
  assign _T_86 = xnor$_io_out_0[15:12];
  assign _T_87 = xnor$_io_out_0[19:16];
  assign _T_88 = xnor$_io_out_0[23:20];
  assign _T_89 = xnor$_io_out_0[27:24];
  assign _T_90 = xnor$_io_out_0[31:28];
  assign _T_141_0 = _T_93;
  assign _T_141_1 = _T_96;
  assign _T_141_2 = _T_99;
  assign _T_141_3 = _T_102;
  assign _T_141_4 = _T_105;
  assign _T_141_5 = _T_108;
  assign _T_141_6 = _T_111;
  assign _T_141_7 = _T_114;
  assign _T_141_8 = _T_117;
  assign _T_141_9 = _T_120;
  assign _T_141_10 = _T_123;
  assign _T_141_11 = _T_126;
  assign _T_141_12 = _T_129;
  assign _T_141_13 = _T_132;
  assign _T_141_14 = _T_135;
  assign _T_141_15 = _T_138;
  assign _T_211_0 = _T_163;
  assign _T_211_1 = _T_166;
  assign _T_211_2 = _T_169;
  assign _T_211_3 = _T_172;
  assign _T_211_4 = _T_175;
  assign _T_211_5 = _T_178;
  assign _T_211_6 = _T_181;
  assign _T_211_7 = _T_184;
  assign _T_211_8 = _T_187;
  assign _T_211_9 = _T_190;
  assign _T_211_10 = _T_193;
  assign _T_211_11 = _T_196;
  assign _T_211_12 = _T_199;
  assign _T_211_13 = _T_202;
  assign _T_211_14 = _T_205;
  assign _T_211_15 = _T_208;
  assign _T_281_0 = _T_233;
  assign _T_281_1 = _T_236;
  assign _T_281_2 = _T_239;
  assign _T_281_3 = _T_242;
  assign _T_281_4 = _T_245;
  assign _T_281_5 = _T_248;
  assign _T_281_6 = _T_251;
  assign _T_281_7 = _T_254;
  assign _T_281_8 = _T_257;
  assign _T_281_9 = _T_260;
  assign _T_281_10 = _T_263;
  assign _T_281_11 = _T_266;
  assign _T_281_12 = _T_269;
  assign _T_281_13 = _T_272;
  assign _T_281_14 = _T_275;
  assign _T_281_15 = _T_278;
  assign _T_351_0 = _T_303;
  assign _T_351_1 = _T_306;
  assign _T_351_2 = _T_309;
  assign _T_351_3 = _T_312;
  assign _T_351_4 = _T_315;
  assign _T_351_5 = _T_318;
  assign _T_351_6 = _T_321;
  assign _T_351_7 = _T_324;
  assign _T_351_8 = _T_327;
  assign _T_351_9 = _T_330;
  assign _T_351_10 = _T_333;
  assign _T_351_11 = _T_336;
  assign _T_351_12 = _T_339;
  assign _T_351_13 = _T_342;
  assign _T_351_14 = _T_345;
  assign _T_351_15 = _T_348;
  assign _T_421_0 = _T_373;
  assign _T_421_1 = _T_376;
  assign _T_421_2 = _T_379;
  assign _T_421_3 = _T_382;
  assign _T_421_4 = _T_385;
  assign _T_421_5 = _T_388;
  assign _T_421_6 = _T_391;
  assign _T_421_7 = _T_394;
  assign _T_421_8 = _T_397;
  assign _T_421_9 = _T_400;
  assign _T_421_10 = _T_403;
  assign _T_421_11 = _T_406;
  assign _T_421_12 = _T_409;
  assign _T_421_13 = _T_412;
  assign _T_421_14 = _T_415;
  assign _T_421_15 = _T_418;
  assign _T_491_0 = _T_443;
  assign _T_491_1 = _T_446;
  assign _T_491_2 = _T_449;
  assign _T_491_3 = _T_452;
  assign _T_491_4 = _T_455;
  assign _T_491_5 = _T_458;
  assign _T_491_6 = _T_461;
  assign _T_491_7 = _T_464;
  assign _T_491_8 = _T_467;
  assign _T_491_9 = _T_470;
  assign _T_491_10 = _T_473;
  assign _T_491_11 = _T_476;
  assign _T_491_12 = _T_479;
  assign _T_491_13 = _T_482;
  assign _T_491_14 = _T_485;
  assign _T_491_15 = _T_488;
  assign _T_561_0 = _T_513;
  assign _T_561_1 = _T_516;
  assign _T_561_2 = _T_519;
  assign _T_561_3 = _T_522;
  assign _T_561_4 = _T_525;
  assign _T_561_5 = _T_528;
  assign _T_561_6 = _T_531;
  assign _T_561_7 = _T_534;
  assign _T_561_8 = _T_537;
  assign _T_561_9 = _T_540;
  assign _T_561_10 = _T_543;
  assign _T_561_11 = _T_546;
  assign _T_561_12 = _T_549;
  assign _T_561_13 = _T_552;
  assign _T_561_14 = _T_555;
  assign _T_561_15 = _T_558;
  assign _T_631_0 = _T_583;
  assign _T_631_1 = _T_586;
  assign _T_631_2 = _T_589;
  assign _T_631_3 = _T_592;
  assign _T_631_4 = _T_595;
  assign _T_631_5 = _T_598;
  assign _T_631_6 = _T_601;
  assign _T_631_7 = _T_604;
  assign _T_631_8 = _T_607;
  assign _T_631_9 = _T_610;
  assign _T_631_10 = _T_613;
  assign _T_631_11 = _T_616;
  assign _T_631_12 = _T_619;
  assign _T_631_13 = _T_622;
  assign _T_631_14 = _T_625;
  assign _T_631_15 = _T_628;
  assign _GEN_0 = _GEN_46;
  assign _GEN_32 = 4'h1 == _T_83 ? $signed(_T_141_1) : $signed(_T_141_0);
  assign _GEN_33 = 4'h2 == _T_83 ? $signed(_T_141_2) : $signed(_GEN_32);
  assign _GEN_34 = 4'h3 == _T_83 ? $signed(_T_141_3) : $signed(_GEN_33);
  assign _GEN_35 = 4'h4 == _T_83 ? $signed(_T_141_4) : $signed(_GEN_34);
  assign _GEN_36 = 4'h5 == _T_83 ? $signed(_T_141_5) : $signed(_GEN_35);
  assign _GEN_37 = 4'h6 == _T_83 ? $signed(_T_141_6) : $signed(_GEN_36);
  assign _GEN_38 = 4'h7 == _T_83 ? $signed(_T_141_7) : $signed(_GEN_37);
  assign _GEN_39 = 4'h8 == _T_83 ? $signed(_T_141_8) : $signed(_GEN_38);
  assign _GEN_40 = 4'h9 == _T_83 ? $signed(_T_141_9) : $signed(_GEN_39);
  assign _GEN_41 = 4'ha == _T_83 ? $signed(_T_141_10) : $signed(_GEN_40);
  assign _GEN_42 = 4'hb == _T_83 ? $signed(_T_141_11) : $signed(_GEN_41);
  assign _GEN_43 = 4'hc == _T_83 ? $signed(_T_141_12) : $signed(_GEN_42);
  assign _GEN_44 = 4'hd == _T_83 ? $signed(_T_141_13) : $signed(_GEN_43);
  assign _GEN_45 = 4'he == _T_83 ? $signed(_T_141_14) : $signed(_GEN_44);
  assign _GEN_46 = 4'hf == _T_83 ? $signed(_T_141_15) : $signed(_GEN_45);
  assign _GEN_1 = _GEN_61;
  assign _GEN_47 = 4'h1 == _T_84 ? $signed(_T_211_1) : $signed(_T_211_0);
  assign _GEN_48 = 4'h2 == _T_84 ? $signed(_T_211_2) : $signed(_GEN_47);
  assign _GEN_49 = 4'h3 == _T_84 ? $signed(_T_211_3) : $signed(_GEN_48);
  assign _GEN_50 = 4'h4 == _T_84 ? $signed(_T_211_4) : $signed(_GEN_49);
  assign _GEN_51 = 4'h5 == _T_84 ? $signed(_T_211_5) : $signed(_GEN_50);
  assign _GEN_52 = 4'h6 == _T_84 ? $signed(_T_211_6) : $signed(_GEN_51);
  assign _GEN_53 = 4'h7 == _T_84 ? $signed(_T_211_7) : $signed(_GEN_52);
  assign _GEN_54 = 4'h8 == _T_84 ? $signed(_T_211_8) : $signed(_GEN_53);
  assign _GEN_55 = 4'h9 == _T_84 ? $signed(_T_211_9) : $signed(_GEN_54);
  assign _GEN_56 = 4'ha == _T_84 ? $signed(_T_211_10) : $signed(_GEN_55);
  assign _GEN_57 = 4'hb == _T_84 ? $signed(_T_211_11) : $signed(_GEN_56);
  assign _GEN_58 = 4'hc == _T_84 ? $signed(_T_211_12) : $signed(_GEN_57);
  assign _GEN_59 = 4'hd == _T_84 ? $signed(_T_211_13) : $signed(_GEN_58);
  assign _GEN_60 = 4'he == _T_84 ? $signed(_T_211_14) : $signed(_GEN_59);
  assign _GEN_61 = 4'hf == _T_84 ? $signed(_T_211_15) : $signed(_GEN_60);
  assign _T_651 = $signed(_GEN_0) + $signed(_GEN_1);
  assign _T_652 = _T_651[5:0];
  assign _T_653 = $signed(_T_652);
  assign _GEN_2 = _GEN_76;
  assign _GEN_62 = 4'h1 == _T_85 ? $signed(_T_281_1) : $signed(_T_281_0);
  assign _GEN_63 = 4'h2 == _T_85 ? $signed(_T_281_2) : $signed(_GEN_62);
  assign _GEN_64 = 4'h3 == _T_85 ? $signed(_T_281_3) : $signed(_GEN_63);
  assign _GEN_65 = 4'h4 == _T_85 ? $signed(_T_281_4) : $signed(_GEN_64);
  assign _GEN_66 = 4'h5 == _T_85 ? $signed(_T_281_5) : $signed(_GEN_65);
  assign _GEN_67 = 4'h6 == _T_85 ? $signed(_T_281_6) : $signed(_GEN_66);
  assign _GEN_68 = 4'h7 == _T_85 ? $signed(_T_281_7) : $signed(_GEN_67);
  assign _GEN_69 = 4'h8 == _T_85 ? $signed(_T_281_8) : $signed(_GEN_68);
  assign _GEN_70 = 4'h9 == _T_85 ? $signed(_T_281_9) : $signed(_GEN_69);
  assign _GEN_71 = 4'ha == _T_85 ? $signed(_T_281_10) : $signed(_GEN_70);
  assign _GEN_72 = 4'hb == _T_85 ? $signed(_T_281_11) : $signed(_GEN_71);
  assign _GEN_73 = 4'hc == _T_85 ? $signed(_T_281_12) : $signed(_GEN_72);
  assign _GEN_74 = 4'hd == _T_85 ? $signed(_T_281_13) : $signed(_GEN_73);
  assign _GEN_75 = 4'he == _T_85 ? $signed(_T_281_14) : $signed(_GEN_74);
  assign _GEN_76 = 4'hf == _T_85 ? $signed(_T_281_15) : $signed(_GEN_75);
  assign _GEN_3 = _GEN_91;
  assign _GEN_77 = 4'h1 == _T_86 ? $signed(_T_351_1) : $signed(_T_351_0);
  assign _GEN_78 = 4'h2 == _T_86 ? $signed(_T_351_2) : $signed(_GEN_77);
  assign _GEN_79 = 4'h3 == _T_86 ? $signed(_T_351_3) : $signed(_GEN_78);
  assign _GEN_80 = 4'h4 == _T_86 ? $signed(_T_351_4) : $signed(_GEN_79);
  assign _GEN_81 = 4'h5 == _T_86 ? $signed(_T_351_5) : $signed(_GEN_80);
  assign _GEN_82 = 4'h6 == _T_86 ? $signed(_T_351_6) : $signed(_GEN_81);
  assign _GEN_83 = 4'h7 == _T_86 ? $signed(_T_351_7) : $signed(_GEN_82);
  assign _GEN_84 = 4'h8 == _T_86 ? $signed(_T_351_8) : $signed(_GEN_83);
  assign _GEN_85 = 4'h9 == _T_86 ? $signed(_T_351_9) : $signed(_GEN_84);
  assign _GEN_86 = 4'ha == _T_86 ? $signed(_T_351_10) : $signed(_GEN_85);
  assign _GEN_87 = 4'hb == _T_86 ? $signed(_T_351_11) : $signed(_GEN_86);
  assign _GEN_88 = 4'hc == _T_86 ? $signed(_T_351_12) : $signed(_GEN_87);
  assign _GEN_89 = 4'hd == _T_86 ? $signed(_T_351_13) : $signed(_GEN_88);
  assign _GEN_90 = 4'he == _T_86 ? $signed(_T_351_14) : $signed(_GEN_89);
  assign _GEN_91 = 4'hf == _T_86 ? $signed(_T_351_15) : $signed(_GEN_90);
  assign _T_654 = $signed(_GEN_2) + $signed(_GEN_3);
  assign _T_655 = _T_654[5:0];
  assign _T_656 = $signed(_T_655);
  assign _GEN_4 = _GEN_106;
  assign _GEN_92 = 4'h1 == _T_87 ? $signed(_T_421_1) : $signed(_T_421_0);
  assign _GEN_93 = 4'h2 == _T_87 ? $signed(_T_421_2) : $signed(_GEN_92);
  assign _GEN_94 = 4'h3 == _T_87 ? $signed(_T_421_3) : $signed(_GEN_93);
  assign _GEN_95 = 4'h4 == _T_87 ? $signed(_T_421_4) : $signed(_GEN_94);
  assign _GEN_96 = 4'h5 == _T_87 ? $signed(_T_421_5) : $signed(_GEN_95);
  assign _GEN_97 = 4'h6 == _T_87 ? $signed(_T_421_6) : $signed(_GEN_96);
  assign _GEN_98 = 4'h7 == _T_87 ? $signed(_T_421_7) : $signed(_GEN_97);
  assign _GEN_99 = 4'h8 == _T_87 ? $signed(_T_421_8) : $signed(_GEN_98);
  assign _GEN_100 = 4'h9 == _T_87 ? $signed(_T_421_9) : $signed(_GEN_99);
  assign _GEN_101 = 4'ha == _T_87 ? $signed(_T_421_10) : $signed(_GEN_100);
  assign _GEN_102 = 4'hb == _T_87 ? $signed(_T_421_11) : $signed(_GEN_101);
  assign _GEN_103 = 4'hc == _T_87 ? $signed(_T_421_12) : $signed(_GEN_102);
  assign _GEN_104 = 4'hd == _T_87 ? $signed(_T_421_13) : $signed(_GEN_103);
  assign _GEN_105 = 4'he == _T_87 ? $signed(_T_421_14) : $signed(_GEN_104);
  assign _GEN_106 = 4'hf == _T_87 ? $signed(_T_421_15) : $signed(_GEN_105);
  assign _GEN_5 = _GEN_121;
  assign _GEN_107 = 4'h1 == _T_88 ? $signed(_T_491_1) : $signed(_T_491_0);
  assign _GEN_108 = 4'h2 == _T_88 ? $signed(_T_491_2) : $signed(_GEN_107);
  assign _GEN_109 = 4'h3 == _T_88 ? $signed(_T_491_3) : $signed(_GEN_108);
  assign _GEN_110 = 4'h4 == _T_88 ? $signed(_T_491_4) : $signed(_GEN_109);
  assign _GEN_111 = 4'h5 == _T_88 ? $signed(_T_491_5) : $signed(_GEN_110);
  assign _GEN_112 = 4'h6 == _T_88 ? $signed(_T_491_6) : $signed(_GEN_111);
  assign _GEN_113 = 4'h7 == _T_88 ? $signed(_T_491_7) : $signed(_GEN_112);
  assign _GEN_114 = 4'h8 == _T_88 ? $signed(_T_491_8) : $signed(_GEN_113);
  assign _GEN_115 = 4'h9 == _T_88 ? $signed(_T_491_9) : $signed(_GEN_114);
  assign _GEN_116 = 4'ha == _T_88 ? $signed(_T_491_10) : $signed(_GEN_115);
  assign _GEN_117 = 4'hb == _T_88 ? $signed(_T_491_11) : $signed(_GEN_116);
  assign _GEN_118 = 4'hc == _T_88 ? $signed(_T_491_12) : $signed(_GEN_117);
  assign _GEN_119 = 4'hd == _T_88 ? $signed(_T_491_13) : $signed(_GEN_118);
  assign _GEN_120 = 4'he == _T_88 ? $signed(_T_491_14) : $signed(_GEN_119);
  assign _GEN_121 = 4'hf == _T_88 ? $signed(_T_491_15) : $signed(_GEN_120);
  assign _T_657 = $signed(_GEN_4) + $signed(_GEN_5);
  assign _T_658 = _T_657[5:0];
  assign _T_659 = $signed(_T_658);
  assign _GEN_6 = _GEN_136;
  assign _GEN_122 = 4'h1 == _T_89 ? $signed(_T_561_1) : $signed(_T_561_0);
  assign _GEN_123 = 4'h2 == _T_89 ? $signed(_T_561_2) : $signed(_GEN_122);
  assign _GEN_124 = 4'h3 == _T_89 ? $signed(_T_561_3) : $signed(_GEN_123);
  assign _GEN_125 = 4'h4 == _T_89 ? $signed(_T_561_4) : $signed(_GEN_124);
  assign _GEN_126 = 4'h5 == _T_89 ? $signed(_T_561_5) : $signed(_GEN_125);
  assign _GEN_127 = 4'h6 == _T_89 ? $signed(_T_561_6) : $signed(_GEN_126);
  assign _GEN_128 = 4'h7 == _T_89 ? $signed(_T_561_7) : $signed(_GEN_127);
  assign _GEN_129 = 4'h8 == _T_89 ? $signed(_T_561_8) : $signed(_GEN_128);
  assign _GEN_130 = 4'h9 == _T_89 ? $signed(_T_561_9) : $signed(_GEN_129);
  assign _GEN_131 = 4'ha == _T_89 ? $signed(_T_561_10) : $signed(_GEN_130);
  assign _GEN_132 = 4'hb == _T_89 ? $signed(_T_561_11) : $signed(_GEN_131);
  assign _GEN_133 = 4'hc == _T_89 ? $signed(_T_561_12) : $signed(_GEN_132);
  assign _GEN_134 = 4'hd == _T_89 ? $signed(_T_561_13) : $signed(_GEN_133);
  assign _GEN_135 = 4'he == _T_89 ? $signed(_T_561_14) : $signed(_GEN_134);
  assign _GEN_136 = 4'hf == _T_89 ? $signed(_T_561_15) : $signed(_GEN_135);
  assign _GEN_7 = _GEN_151;
  assign _GEN_137 = 4'h1 == _T_90 ? $signed(_T_631_1) : $signed(_T_631_0);
  assign _GEN_138 = 4'h2 == _T_90 ? $signed(_T_631_2) : $signed(_GEN_137);
  assign _GEN_139 = 4'h3 == _T_90 ? $signed(_T_631_3) : $signed(_GEN_138);
  assign _GEN_140 = 4'h4 == _T_90 ? $signed(_T_631_4) : $signed(_GEN_139);
  assign _GEN_141 = 4'h5 == _T_90 ? $signed(_T_631_5) : $signed(_GEN_140);
  assign _GEN_142 = 4'h6 == _T_90 ? $signed(_T_631_6) : $signed(_GEN_141);
  assign _GEN_143 = 4'h7 == _T_90 ? $signed(_T_631_7) : $signed(_GEN_142);
  assign _GEN_144 = 4'h8 == _T_90 ? $signed(_T_631_8) : $signed(_GEN_143);
  assign _GEN_145 = 4'h9 == _T_90 ? $signed(_T_631_9) : $signed(_GEN_144);
  assign _GEN_146 = 4'ha == _T_90 ? $signed(_T_631_10) : $signed(_GEN_145);
  assign _GEN_147 = 4'hb == _T_90 ? $signed(_T_631_11) : $signed(_GEN_146);
  assign _GEN_148 = 4'hc == _T_90 ? $signed(_T_631_12) : $signed(_GEN_147);
  assign _GEN_149 = 4'hd == _T_90 ? $signed(_T_631_13) : $signed(_GEN_148);
  assign _GEN_150 = 4'he == _T_90 ? $signed(_T_631_14) : $signed(_GEN_149);
  assign _GEN_151 = 4'hf == _T_90 ? $signed(_T_631_15) : $signed(_GEN_150);
  assign _T_660 = $signed(_GEN_6) + $signed(_GEN_7);
  assign _T_661 = _T_660[5:0];
  assign _T_662 = $signed(_T_661);
  assign _T_663 = $signed(_T_653) + $signed(_T_656);
  assign _T_664 = _T_663[5:0];
  assign _T_665 = $signed(_T_664);
  assign _T_666 = $signed(_T_659) + $signed(_T_662);
  assign _T_667 = _T_666[5:0];
  assign _T_668 = $signed(_T_667);
  assign _T_669 = $signed(_T_665) + $signed(_T_668);
  assign _T_670 = _T_669[5:0];
  assign _T_671 = $signed(_T_670);
  assign MulAdd_io_a = _T_676;
  assign MulAdd_io_b = $signed(_GEN_512);
  assign MulAdd_io_m = mean_io_output;
  assign MulAdd_io_c = _T_678;
  assign _T_673 = mem_io_out[127:96];
  assign _T_674 = io_memSel ? 32'h0 : _T_673;
  assign _T_675 = _T_674[31:16];
  assign _T_676 = $signed(_T_675);
  assign _T_677 = _T_674[15:0];
  assign _T_678 = $signed(_T_677);
  assign signs_0 = MulAdd_io_r[31];
  assign Accumulator_1_clock = clock;
  assign Accumulator_1_io_in = {{26{_T_1267[5]}},_T_1267};
  assign Accumulator_1_io_sel = io_accSel;
  assign Accumulator_1_io_en = io_accEn;
  assign Accumulator_1_io_reset = io_accReset;
  assign _T_679 = xnor$_io_out_1[3:0];
  assign _T_680 = xnor$_io_out_1[7:4];
  assign _T_681 = xnor$_io_out_1[11:8];
  assign _T_682 = xnor$_io_out_1[15:12];
  assign _T_683 = xnor$_io_out_1[19:16];
  assign _T_684 = xnor$_io_out_1[23:20];
  assign _T_685 = xnor$_io_out_1[27:24];
  assign _T_686 = xnor$_io_out_1[31:28];
  assign _T_737_0 = _T_689;
  assign _T_737_1 = _T_692;
  assign _T_737_2 = _T_695;
  assign _T_737_3 = _T_698;
  assign _T_737_4 = _T_701;
  assign _T_737_5 = _T_704;
  assign _T_737_6 = _T_707;
  assign _T_737_7 = _T_710;
  assign _T_737_8 = _T_713;
  assign _T_737_9 = _T_716;
  assign _T_737_10 = _T_719;
  assign _T_737_11 = _T_722;
  assign _T_737_12 = _T_725;
  assign _T_737_13 = _T_728;
  assign _T_737_14 = _T_731;
  assign _T_737_15 = _T_734;
  assign _T_807_0 = _T_759;
  assign _T_807_1 = _T_762;
  assign _T_807_2 = _T_765;
  assign _T_807_3 = _T_768;
  assign _T_807_4 = _T_771;
  assign _T_807_5 = _T_774;
  assign _T_807_6 = _T_777;
  assign _T_807_7 = _T_780;
  assign _T_807_8 = _T_783;
  assign _T_807_9 = _T_786;
  assign _T_807_10 = _T_789;
  assign _T_807_11 = _T_792;
  assign _T_807_12 = _T_795;
  assign _T_807_13 = _T_798;
  assign _T_807_14 = _T_801;
  assign _T_807_15 = _T_804;
  assign _T_877_0 = _T_829;
  assign _T_877_1 = _T_832;
  assign _T_877_2 = _T_835;
  assign _T_877_3 = _T_838;
  assign _T_877_4 = _T_841;
  assign _T_877_5 = _T_844;
  assign _T_877_6 = _T_847;
  assign _T_877_7 = _T_850;
  assign _T_877_8 = _T_853;
  assign _T_877_9 = _T_856;
  assign _T_877_10 = _T_859;
  assign _T_877_11 = _T_862;
  assign _T_877_12 = _T_865;
  assign _T_877_13 = _T_868;
  assign _T_877_14 = _T_871;
  assign _T_877_15 = _T_874;
  assign _T_947_0 = _T_899;
  assign _T_947_1 = _T_902;
  assign _T_947_2 = _T_905;
  assign _T_947_3 = _T_908;
  assign _T_947_4 = _T_911;
  assign _T_947_5 = _T_914;
  assign _T_947_6 = _T_917;
  assign _T_947_7 = _T_920;
  assign _T_947_8 = _T_923;
  assign _T_947_9 = _T_926;
  assign _T_947_10 = _T_929;
  assign _T_947_11 = _T_932;
  assign _T_947_12 = _T_935;
  assign _T_947_13 = _T_938;
  assign _T_947_14 = _T_941;
  assign _T_947_15 = _T_944;
  assign _T_1017_0 = _T_969;
  assign _T_1017_1 = _T_972;
  assign _T_1017_2 = _T_975;
  assign _T_1017_3 = _T_978;
  assign _T_1017_4 = _T_981;
  assign _T_1017_5 = _T_984;
  assign _T_1017_6 = _T_987;
  assign _T_1017_7 = _T_990;
  assign _T_1017_8 = _T_993;
  assign _T_1017_9 = _T_996;
  assign _T_1017_10 = _T_999;
  assign _T_1017_11 = _T_1002;
  assign _T_1017_12 = _T_1005;
  assign _T_1017_13 = _T_1008;
  assign _T_1017_14 = _T_1011;
  assign _T_1017_15 = _T_1014;
  assign _T_1087_0 = _T_1039;
  assign _T_1087_1 = _T_1042;
  assign _T_1087_2 = _T_1045;
  assign _T_1087_3 = _T_1048;
  assign _T_1087_4 = _T_1051;
  assign _T_1087_5 = _T_1054;
  assign _T_1087_6 = _T_1057;
  assign _T_1087_7 = _T_1060;
  assign _T_1087_8 = _T_1063;
  assign _T_1087_9 = _T_1066;
  assign _T_1087_10 = _T_1069;
  assign _T_1087_11 = _T_1072;
  assign _T_1087_12 = _T_1075;
  assign _T_1087_13 = _T_1078;
  assign _T_1087_14 = _T_1081;
  assign _T_1087_15 = _T_1084;
  assign _T_1157_0 = _T_1109;
  assign _T_1157_1 = _T_1112;
  assign _T_1157_2 = _T_1115;
  assign _T_1157_3 = _T_1118;
  assign _T_1157_4 = _T_1121;
  assign _T_1157_5 = _T_1124;
  assign _T_1157_6 = _T_1127;
  assign _T_1157_7 = _T_1130;
  assign _T_1157_8 = _T_1133;
  assign _T_1157_9 = _T_1136;
  assign _T_1157_10 = _T_1139;
  assign _T_1157_11 = _T_1142;
  assign _T_1157_12 = _T_1145;
  assign _T_1157_13 = _T_1148;
  assign _T_1157_14 = _T_1151;
  assign _T_1157_15 = _T_1154;
  assign _T_1227_0 = _T_1179;
  assign _T_1227_1 = _T_1182;
  assign _T_1227_2 = _T_1185;
  assign _T_1227_3 = _T_1188;
  assign _T_1227_4 = _T_1191;
  assign _T_1227_5 = _T_1194;
  assign _T_1227_6 = _T_1197;
  assign _T_1227_7 = _T_1200;
  assign _T_1227_8 = _T_1203;
  assign _T_1227_9 = _T_1206;
  assign _T_1227_10 = _T_1209;
  assign _T_1227_11 = _T_1212;
  assign _T_1227_12 = _T_1215;
  assign _T_1227_13 = _T_1218;
  assign _T_1227_14 = _T_1221;
  assign _T_1227_15 = _T_1224;
  assign _GEN_8 = _GEN_166;
  assign _GEN_152 = 4'h1 == _T_679 ? $signed(_T_737_1) : $signed(_T_737_0);
  assign _GEN_153 = 4'h2 == _T_679 ? $signed(_T_737_2) : $signed(_GEN_152);
  assign _GEN_154 = 4'h3 == _T_679 ? $signed(_T_737_3) : $signed(_GEN_153);
  assign _GEN_155 = 4'h4 == _T_679 ? $signed(_T_737_4) : $signed(_GEN_154);
  assign _GEN_156 = 4'h5 == _T_679 ? $signed(_T_737_5) : $signed(_GEN_155);
  assign _GEN_157 = 4'h6 == _T_679 ? $signed(_T_737_6) : $signed(_GEN_156);
  assign _GEN_158 = 4'h7 == _T_679 ? $signed(_T_737_7) : $signed(_GEN_157);
  assign _GEN_159 = 4'h8 == _T_679 ? $signed(_T_737_8) : $signed(_GEN_158);
  assign _GEN_160 = 4'h9 == _T_679 ? $signed(_T_737_9) : $signed(_GEN_159);
  assign _GEN_161 = 4'ha == _T_679 ? $signed(_T_737_10) : $signed(_GEN_160);
  assign _GEN_162 = 4'hb == _T_679 ? $signed(_T_737_11) : $signed(_GEN_161);
  assign _GEN_163 = 4'hc == _T_679 ? $signed(_T_737_12) : $signed(_GEN_162);
  assign _GEN_164 = 4'hd == _T_679 ? $signed(_T_737_13) : $signed(_GEN_163);
  assign _GEN_165 = 4'he == _T_679 ? $signed(_T_737_14) : $signed(_GEN_164);
  assign _GEN_166 = 4'hf == _T_679 ? $signed(_T_737_15) : $signed(_GEN_165);
  assign _GEN_9 = _GEN_181;
  assign _GEN_167 = 4'h1 == _T_680 ? $signed(_T_807_1) : $signed(_T_807_0);
  assign _GEN_168 = 4'h2 == _T_680 ? $signed(_T_807_2) : $signed(_GEN_167);
  assign _GEN_169 = 4'h3 == _T_680 ? $signed(_T_807_3) : $signed(_GEN_168);
  assign _GEN_170 = 4'h4 == _T_680 ? $signed(_T_807_4) : $signed(_GEN_169);
  assign _GEN_171 = 4'h5 == _T_680 ? $signed(_T_807_5) : $signed(_GEN_170);
  assign _GEN_172 = 4'h6 == _T_680 ? $signed(_T_807_6) : $signed(_GEN_171);
  assign _GEN_173 = 4'h7 == _T_680 ? $signed(_T_807_7) : $signed(_GEN_172);
  assign _GEN_174 = 4'h8 == _T_680 ? $signed(_T_807_8) : $signed(_GEN_173);
  assign _GEN_175 = 4'h9 == _T_680 ? $signed(_T_807_9) : $signed(_GEN_174);
  assign _GEN_176 = 4'ha == _T_680 ? $signed(_T_807_10) : $signed(_GEN_175);
  assign _GEN_177 = 4'hb == _T_680 ? $signed(_T_807_11) : $signed(_GEN_176);
  assign _GEN_178 = 4'hc == _T_680 ? $signed(_T_807_12) : $signed(_GEN_177);
  assign _GEN_179 = 4'hd == _T_680 ? $signed(_T_807_13) : $signed(_GEN_178);
  assign _GEN_180 = 4'he == _T_680 ? $signed(_T_807_14) : $signed(_GEN_179);
  assign _GEN_181 = 4'hf == _T_680 ? $signed(_T_807_15) : $signed(_GEN_180);
  assign _T_1247 = $signed(_GEN_8) + $signed(_GEN_9);
  assign _T_1248 = _T_1247[5:0];
  assign _T_1249 = $signed(_T_1248);
  assign _GEN_10 = _GEN_196;
  assign _GEN_182 = 4'h1 == _T_681 ? $signed(_T_877_1) : $signed(_T_877_0);
  assign _GEN_183 = 4'h2 == _T_681 ? $signed(_T_877_2) : $signed(_GEN_182);
  assign _GEN_184 = 4'h3 == _T_681 ? $signed(_T_877_3) : $signed(_GEN_183);
  assign _GEN_185 = 4'h4 == _T_681 ? $signed(_T_877_4) : $signed(_GEN_184);
  assign _GEN_186 = 4'h5 == _T_681 ? $signed(_T_877_5) : $signed(_GEN_185);
  assign _GEN_187 = 4'h6 == _T_681 ? $signed(_T_877_6) : $signed(_GEN_186);
  assign _GEN_188 = 4'h7 == _T_681 ? $signed(_T_877_7) : $signed(_GEN_187);
  assign _GEN_189 = 4'h8 == _T_681 ? $signed(_T_877_8) : $signed(_GEN_188);
  assign _GEN_190 = 4'h9 == _T_681 ? $signed(_T_877_9) : $signed(_GEN_189);
  assign _GEN_191 = 4'ha == _T_681 ? $signed(_T_877_10) : $signed(_GEN_190);
  assign _GEN_192 = 4'hb == _T_681 ? $signed(_T_877_11) : $signed(_GEN_191);
  assign _GEN_193 = 4'hc == _T_681 ? $signed(_T_877_12) : $signed(_GEN_192);
  assign _GEN_194 = 4'hd == _T_681 ? $signed(_T_877_13) : $signed(_GEN_193);
  assign _GEN_195 = 4'he == _T_681 ? $signed(_T_877_14) : $signed(_GEN_194);
  assign _GEN_196 = 4'hf == _T_681 ? $signed(_T_877_15) : $signed(_GEN_195);
  assign _GEN_11 = _GEN_211;
  assign _GEN_197 = 4'h1 == _T_682 ? $signed(_T_947_1) : $signed(_T_947_0);
  assign _GEN_198 = 4'h2 == _T_682 ? $signed(_T_947_2) : $signed(_GEN_197);
  assign _GEN_199 = 4'h3 == _T_682 ? $signed(_T_947_3) : $signed(_GEN_198);
  assign _GEN_200 = 4'h4 == _T_682 ? $signed(_T_947_4) : $signed(_GEN_199);
  assign _GEN_201 = 4'h5 == _T_682 ? $signed(_T_947_5) : $signed(_GEN_200);
  assign _GEN_202 = 4'h6 == _T_682 ? $signed(_T_947_6) : $signed(_GEN_201);
  assign _GEN_203 = 4'h7 == _T_682 ? $signed(_T_947_7) : $signed(_GEN_202);
  assign _GEN_204 = 4'h8 == _T_682 ? $signed(_T_947_8) : $signed(_GEN_203);
  assign _GEN_205 = 4'h9 == _T_682 ? $signed(_T_947_9) : $signed(_GEN_204);
  assign _GEN_206 = 4'ha == _T_682 ? $signed(_T_947_10) : $signed(_GEN_205);
  assign _GEN_207 = 4'hb == _T_682 ? $signed(_T_947_11) : $signed(_GEN_206);
  assign _GEN_208 = 4'hc == _T_682 ? $signed(_T_947_12) : $signed(_GEN_207);
  assign _GEN_209 = 4'hd == _T_682 ? $signed(_T_947_13) : $signed(_GEN_208);
  assign _GEN_210 = 4'he == _T_682 ? $signed(_T_947_14) : $signed(_GEN_209);
  assign _GEN_211 = 4'hf == _T_682 ? $signed(_T_947_15) : $signed(_GEN_210);
  assign _T_1250 = $signed(_GEN_10) + $signed(_GEN_11);
  assign _T_1251 = _T_1250[5:0];
  assign _T_1252 = $signed(_T_1251);
  assign _GEN_12 = _GEN_226;
  assign _GEN_212 = 4'h1 == _T_683 ? $signed(_T_1017_1) : $signed(_T_1017_0);
  assign _GEN_213 = 4'h2 == _T_683 ? $signed(_T_1017_2) : $signed(_GEN_212);
  assign _GEN_214 = 4'h3 == _T_683 ? $signed(_T_1017_3) : $signed(_GEN_213);
  assign _GEN_215 = 4'h4 == _T_683 ? $signed(_T_1017_4) : $signed(_GEN_214);
  assign _GEN_216 = 4'h5 == _T_683 ? $signed(_T_1017_5) : $signed(_GEN_215);
  assign _GEN_217 = 4'h6 == _T_683 ? $signed(_T_1017_6) : $signed(_GEN_216);
  assign _GEN_218 = 4'h7 == _T_683 ? $signed(_T_1017_7) : $signed(_GEN_217);
  assign _GEN_219 = 4'h8 == _T_683 ? $signed(_T_1017_8) : $signed(_GEN_218);
  assign _GEN_220 = 4'h9 == _T_683 ? $signed(_T_1017_9) : $signed(_GEN_219);
  assign _GEN_221 = 4'ha == _T_683 ? $signed(_T_1017_10) : $signed(_GEN_220);
  assign _GEN_222 = 4'hb == _T_683 ? $signed(_T_1017_11) : $signed(_GEN_221);
  assign _GEN_223 = 4'hc == _T_683 ? $signed(_T_1017_12) : $signed(_GEN_222);
  assign _GEN_224 = 4'hd == _T_683 ? $signed(_T_1017_13) : $signed(_GEN_223);
  assign _GEN_225 = 4'he == _T_683 ? $signed(_T_1017_14) : $signed(_GEN_224);
  assign _GEN_226 = 4'hf == _T_683 ? $signed(_T_1017_15) : $signed(_GEN_225);
  assign _GEN_13 = _GEN_241;
  assign _GEN_227 = 4'h1 == _T_684 ? $signed(_T_1087_1) : $signed(_T_1087_0);
  assign _GEN_228 = 4'h2 == _T_684 ? $signed(_T_1087_2) : $signed(_GEN_227);
  assign _GEN_229 = 4'h3 == _T_684 ? $signed(_T_1087_3) : $signed(_GEN_228);
  assign _GEN_230 = 4'h4 == _T_684 ? $signed(_T_1087_4) : $signed(_GEN_229);
  assign _GEN_231 = 4'h5 == _T_684 ? $signed(_T_1087_5) : $signed(_GEN_230);
  assign _GEN_232 = 4'h6 == _T_684 ? $signed(_T_1087_6) : $signed(_GEN_231);
  assign _GEN_233 = 4'h7 == _T_684 ? $signed(_T_1087_7) : $signed(_GEN_232);
  assign _GEN_234 = 4'h8 == _T_684 ? $signed(_T_1087_8) : $signed(_GEN_233);
  assign _GEN_235 = 4'h9 == _T_684 ? $signed(_T_1087_9) : $signed(_GEN_234);
  assign _GEN_236 = 4'ha == _T_684 ? $signed(_T_1087_10) : $signed(_GEN_235);
  assign _GEN_237 = 4'hb == _T_684 ? $signed(_T_1087_11) : $signed(_GEN_236);
  assign _GEN_238 = 4'hc == _T_684 ? $signed(_T_1087_12) : $signed(_GEN_237);
  assign _GEN_239 = 4'hd == _T_684 ? $signed(_T_1087_13) : $signed(_GEN_238);
  assign _GEN_240 = 4'he == _T_684 ? $signed(_T_1087_14) : $signed(_GEN_239);
  assign _GEN_241 = 4'hf == _T_684 ? $signed(_T_1087_15) : $signed(_GEN_240);
  assign _T_1253 = $signed(_GEN_12) + $signed(_GEN_13);
  assign _T_1254 = _T_1253[5:0];
  assign _T_1255 = $signed(_T_1254);
  assign _GEN_14 = _GEN_256;
  assign _GEN_242 = 4'h1 == _T_685 ? $signed(_T_1157_1) : $signed(_T_1157_0);
  assign _GEN_243 = 4'h2 == _T_685 ? $signed(_T_1157_2) : $signed(_GEN_242);
  assign _GEN_244 = 4'h3 == _T_685 ? $signed(_T_1157_3) : $signed(_GEN_243);
  assign _GEN_245 = 4'h4 == _T_685 ? $signed(_T_1157_4) : $signed(_GEN_244);
  assign _GEN_246 = 4'h5 == _T_685 ? $signed(_T_1157_5) : $signed(_GEN_245);
  assign _GEN_247 = 4'h6 == _T_685 ? $signed(_T_1157_6) : $signed(_GEN_246);
  assign _GEN_248 = 4'h7 == _T_685 ? $signed(_T_1157_7) : $signed(_GEN_247);
  assign _GEN_249 = 4'h8 == _T_685 ? $signed(_T_1157_8) : $signed(_GEN_248);
  assign _GEN_250 = 4'h9 == _T_685 ? $signed(_T_1157_9) : $signed(_GEN_249);
  assign _GEN_251 = 4'ha == _T_685 ? $signed(_T_1157_10) : $signed(_GEN_250);
  assign _GEN_252 = 4'hb == _T_685 ? $signed(_T_1157_11) : $signed(_GEN_251);
  assign _GEN_253 = 4'hc == _T_685 ? $signed(_T_1157_12) : $signed(_GEN_252);
  assign _GEN_254 = 4'hd == _T_685 ? $signed(_T_1157_13) : $signed(_GEN_253);
  assign _GEN_255 = 4'he == _T_685 ? $signed(_T_1157_14) : $signed(_GEN_254);
  assign _GEN_256 = 4'hf == _T_685 ? $signed(_T_1157_15) : $signed(_GEN_255);
  assign _GEN_15 = _GEN_271;
  assign _GEN_257 = 4'h1 == _T_686 ? $signed(_T_1227_1) : $signed(_T_1227_0);
  assign _GEN_258 = 4'h2 == _T_686 ? $signed(_T_1227_2) : $signed(_GEN_257);
  assign _GEN_259 = 4'h3 == _T_686 ? $signed(_T_1227_3) : $signed(_GEN_258);
  assign _GEN_260 = 4'h4 == _T_686 ? $signed(_T_1227_4) : $signed(_GEN_259);
  assign _GEN_261 = 4'h5 == _T_686 ? $signed(_T_1227_5) : $signed(_GEN_260);
  assign _GEN_262 = 4'h6 == _T_686 ? $signed(_T_1227_6) : $signed(_GEN_261);
  assign _GEN_263 = 4'h7 == _T_686 ? $signed(_T_1227_7) : $signed(_GEN_262);
  assign _GEN_264 = 4'h8 == _T_686 ? $signed(_T_1227_8) : $signed(_GEN_263);
  assign _GEN_265 = 4'h9 == _T_686 ? $signed(_T_1227_9) : $signed(_GEN_264);
  assign _GEN_266 = 4'ha == _T_686 ? $signed(_T_1227_10) : $signed(_GEN_265);
  assign _GEN_267 = 4'hb == _T_686 ? $signed(_T_1227_11) : $signed(_GEN_266);
  assign _GEN_268 = 4'hc == _T_686 ? $signed(_T_1227_12) : $signed(_GEN_267);
  assign _GEN_269 = 4'hd == _T_686 ? $signed(_T_1227_13) : $signed(_GEN_268);
  assign _GEN_270 = 4'he == _T_686 ? $signed(_T_1227_14) : $signed(_GEN_269);
  assign _GEN_271 = 4'hf == _T_686 ? $signed(_T_1227_15) : $signed(_GEN_270);
  assign _T_1256 = $signed(_GEN_14) + $signed(_GEN_15);
  assign _T_1257 = _T_1256[5:0];
  assign _T_1258 = $signed(_T_1257);
  assign _T_1259 = $signed(_T_1249) + $signed(_T_1252);
  assign _T_1260 = _T_1259[5:0];
  assign _T_1261 = $signed(_T_1260);
  assign _T_1262 = $signed(_T_1255) + $signed(_T_1258);
  assign _T_1263 = _T_1262[5:0];
  assign _T_1264 = $signed(_T_1263);
  assign _T_1265 = $signed(_T_1261) + $signed(_T_1264);
  assign _T_1266 = _T_1265[5:0];
  assign _T_1267 = $signed(_T_1266);
  assign MulAdd_1_io_a = _T_1272;
  assign MulAdd_1_io_b = $signed(_GEN_513);
  assign MulAdd_1_io_m = mean_io_output;
  assign MulAdd_1_io_c = _T_1274;
  assign _T_1269 = mem_io_out[95:64];
  assign _T_1270 = io_memSel ? 32'h0 : _T_1269;
  assign _T_1271 = _T_1270[31:16];
  assign _T_1272 = $signed(_T_1271);
  assign _T_1273 = _T_1270[15:0];
  assign _T_1274 = $signed(_T_1273);
  assign signs_1 = MulAdd_1_io_r[31];
  assign Accumulator_2_clock = clock;
  assign Accumulator_2_io_in = {{26{_T_1863[5]}},_T_1863};
  assign Accumulator_2_io_sel = io_accSel;
  assign Accumulator_2_io_en = io_accEn;
  assign Accumulator_2_io_reset = io_accReset;
  assign _T_1275 = xnor$_io_out_2[3:0];
  assign _T_1276 = xnor$_io_out_2[7:4];
  assign _T_1277 = xnor$_io_out_2[11:8];
  assign _T_1278 = xnor$_io_out_2[15:12];
  assign _T_1279 = xnor$_io_out_2[19:16];
  assign _T_1280 = xnor$_io_out_2[23:20];
  assign _T_1281 = xnor$_io_out_2[27:24];
  assign _T_1282 = xnor$_io_out_2[31:28];
  assign _T_1333_0 = _T_1285;
  assign _T_1333_1 = _T_1288;
  assign _T_1333_2 = _T_1291;
  assign _T_1333_3 = _T_1294;
  assign _T_1333_4 = _T_1297;
  assign _T_1333_5 = _T_1300;
  assign _T_1333_6 = _T_1303;
  assign _T_1333_7 = _T_1306;
  assign _T_1333_8 = _T_1309;
  assign _T_1333_9 = _T_1312;
  assign _T_1333_10 = _T_1315;
  assign _T_1333_11 = _T_1318;
  assign _T_1333_12 = _T_1321;
  assign _T_1333_13 = _T_1324;
  assign _T_1333_14 = _T_1327;
  assign _T_1333_15 = _T_1330;
  assign _T_1403_0 = _T_1355;
  assign _T_1403_1 = _T_1358;
  assign _T_1403_2 = _T_1361;
  assign _T_1403_3 = _T_1364;
  assign _T_1403_4 = _T_1367;
  assign _T_1403_5 = _T_1370;
  assign _T_1403_6 = _T_1373;
  assign _T_1403_7 = _T_1376;
  assign _T_1403_8 = _T_1379;
  assign _T_1403_9 = _T_1382;
  assign _T_1403_10 = _T_1385;
  assign _T_1403_11 = _T_1388;
  assign _T_1403_12 = _T_1391;
  assign _T_1403_13 = _T_1394;
  assign _T_1403_14 = _T_1397;
  assign _T_1403_15 = _T_1400;
  assign _T_1473_0 = _T_1425;
  assign _T_1473_1 = _T_1428;
  assign _T_1473_2 = _T_1431;
  assign _T_1473_3 = _T_1434;
  assign _T_1473_4 = _T_1437;
  assign _T_1473_5 = _T_1440;
  assign _T_1473_6 = _T_1443;
  assign _T_1473_7 = _T_1446;
  assign _T_1473_8 = _T_1449;
  assign _T_1473_9 = _T_1452;
  assign _T_1473_10 = _T_1455;
  assign _T_1473_11 = _T_1458;
  assign _T_1473_12 = _T_1461;
  assign _T_1473_13 = _T_1464;
  assign _T_1473_14 = _T_1467;
  assign _T_1473_15 = _T_1470;
  assign _T_1543_0 = _T_1495;
  assign _T_1543_1 = _T_1498;
  assign _T_1543_2 = _T_1501;
  assign _T_1543_3 = _T_1504;
  assign _T_1543_4 = _T_1507;
  assign _T_1543_5 = _T_1510;
  assign _T_1543_6 = _T_1513;
  assign _T_1543_7 = _T_1516;
  assign _T_1543_8 = _T_1519;
  assign _T_1543_9 = _T_1522;
  assign _T_1543_10 = _T_1525;
  assign _T_1543_11 = _T_1528;
  assign _T_1543_12 = _T_1531;
  assign _T_1543_13 = _T_1534;
  assign _T_1543_14 = _T_1537;
  assign _T_1543_15 = _T_1540;
  assign _T_1613_0 = _T_1565;
  assign _T_1613_1 = _T_1568;
  assign _T_1613_2 = _T_1571;
  assign _T_1613_3 = _T_1574;
  assign _T_1613_4 = _T_1577;
  assign _T_1613_5 = _T_1580;
  assign _T_1613_6 = _T_1583;
  assign _T_1613_7 = _T_1586;
  assign _T_1613_8 = _T_1589;
  assign _T_1613_9 = _T_1592;
  assign _T_1613_10 = _T_1595;
  assign _T_1613_11 = _T_1598;
  assign _T_1613_12 = _T_1601;
  assign _T_1613_13 = _T_1604;
  assign _T_1613_14 = _T_1607;
  assign _T_1613_15 = _T_1610;
  assign _T_1683_0 = _T_1635;
  assign _T_1683_1 = _T_1638;
  assign _T_1683_2 = _T_1641;
  assign _T_1683_3 = _T_1644;
  assign _T_1683_4 = _T_1647;
  assign _T_1683_5 = _T_1650;
  assign _T_1683_6 = _T_1653;
  assign _T_1683_7 = _T_1656;
  assign _T_1683_8 = _T_1659;
  assign _T_1683_9 = _T_1662;
  assign _T_1683_10 = _T_1665;
  assign _T_1683_11 = _T_1668;
  assign _T_1683_12 = _T_1671;
  assign _T_1683_13 = _T_1674;
  assign _T_1683_14 = _T_1677;
  assign _T_1683_15 = _T_1680;
  assign _T_1753_0 = _T_1705;
  assign _T_1753_1 = _T_1708;
  assign _T_1753_2 = _T_1711;
  assign _T_1753_3 = _T_1714;
  assign _T_1753_4 = _T_1717;
  assign _T_1753_5 = _T_1720;
  assign _T_1753_6 = _T_1723;
  assign _T_1753_7 = _T_1726;
  assign _T_1753_8 = _T_1729;
  assign _T_1753_9 = _T_1732;
  assign _T_1753_10 = _T_1735;
  assign _T_1753_11 = _T_1738;
  assign _T_1753_12 = _T_1741;
  assign _T_1753_13 = _T_1744;
  assign _T_1753_14 = _T_1747;
  assign _T_1753_15 = _T_1750;
  assign _T_1823_0 = _T_1775;
  assign _T_1823_1 = _T_1778;
  assign _T_1823_2 = _T_1781;
  assign _T_1823_3 = _T_1784;
  assign _T_1823_4 = _T_1787;
  assign _T_1823_5 = _T_1790;
  assign _T_1823_6 = _T_1793;
  assign _T_1823_7 = _T_1796;
  assign _T_1823_8 = _T_1799;
  assign _T_1823_9 = _T_1802;
  assign _T_1823_10 = _T_1805;
  assign _T_1823_11 = _T_1808;
  assign _T_1823_12 = _T_1811;
  assign _T_1823_13 = _T_1814;
  assign _T_1823_14 = _T_1817;
  assign _T_1823_15 = _T_1820;
  assign _GEN_16 = _GEN_286;
  assign _GEN_272 = 4'h1 == _T_1275 ? $signed(_T_1333_1) : $signed(_T_1333_0);
  assign _GEN_273 = 4'h2 == _T_1275 ? $signed(_T_1333_2) : $signed(_GEN_272);
  assign _GEN_274 = 4'h3 == _T_1275 ? $signed(_T_1333_3) : $signed(_GEN_273);
  assign _GEN_275 = 4'h4 == _T_1275 ? $signed(_T_1333_4) : $signed(_GEN_274);
  assign _GEN_276 = 4'h5 == _T_1275 ? $signed(_T_1333_5) : $signed(_GEN_275);
  assign _GEN_277 = 4'h6 == _T_1275 ? $signed(_T_1333_6) : $signed(_GEN_276);
  assign _GEN_278 = 4'h7 == _T_1275 ? $signed(_T_1333_7) : $signed(_GEN_277);
  assign _GEN_279 = 4'h8 == _T_1275 ? $signed(_T_1333_8) : $signed(_GEN_278);
  assign _GEN_280 = 4'h9 == _T_1275 ? $signed(_T_1333_9) : $signed(_GEN_279);
  assign _GEN_281 = 4'ha == _T_1275 ? $signed(_T_1333_10) : $signed(_GEN_280);
  assign _GEN_282 = 4'hb == _T_1275 ? $signed(_T_1333_11) : $signed(_GEN_281);
  assign _GEN_283 = 4'hc == _T_1275 ? $signed(_T_1333_12) : $signed(_GEN_282);
  assign _GEN_284 = 4'hd == _T_1275 ? $signed(_T_1333_13) : $signed(_GEN_283);
  assign _GEN_285 = 4'he == _T_1275 ? $signed(_T_1333_14) : $signed(_GEN_284);
  assign _GEN_286 = 4'hf == _T_1275 ? $signed(_T_1333_15) : $signed(_GEN_285);
  assign _GEN_17 = _GEN_301;
  assign _GEN_287 = 4'h1 == _T_1276 ? $signed(_T_1403_1) : $signed(_T_1403_0);
  assign _GEN_288 = 4'h2 == _T_1276 ? $signed(_T_1403_2) : $signed(_GEN_287);
  assign _GEN_289 = 4'h3 == _T_1276 ? $signed(_T_1403_3) : $signed(_GEN_288);
  assign _GEN_290 = 4'h4 == _T_1276 ? $signed(_T_1403_4) : $signed(_GEN_289);
  assign _GEN_291 = 4'h5 == _T_1276 ? $signed(_T_1403_5) : $signed(_GEN_290);
  assign _GEN_292 = 4'h6 == _T_1276 ? $signed(_T_1403_6) : $signed(_GEN_291);
  assign _GEN_293 = 4'h7 == _T_1276 ? $signed(_T_1403_7) : $signed(_GEN_292);
  assign _GEN_294 = 4'h8 == _T_1276 ? $signed(_T_1403_8) : $signed(_GEN_293);
  assign _GEN_295 = 4'h9 == _T_1276 ? $signed(_T_1403_9) : $signed(_GEN_294);
  assign _GEN_296 = 4'ha == _T_1276 ? $signed(_T_1403_10) : $signed(_GEN_295);
  assign _GEN_297 = 4'hb == _T_1276 ? $signed(_T_1403_11) : $signed(_GEN_296);
  assign _GEN_298 = 4'hc == _T_1276 ? $signed(_T_1403_12) : $signed(_GEN_297);
  assign _GEN_299 = 4'hd == _T_1276 ? $signed(_T_1403_13) : $signed(_GEN_298);
  assign _GEN_300 = 4'he == _T_1276 ? $signed(_T_1403_14) : $signed(_GEN_299);
  assign _GEN_301 = 4'hf == _T_1276 ? $signed(_T_1403_15) : $signed(_GEN_300);
  assign _T_1843 = $signed(_GEN_16) + $signed(_GEN_17);
  assign _T_1844 = _T_1843[5:0];
  assign _T_1845 = $signed(_T_1844);
  assign _GEN_18 = _GEN_316;
  assign _GEN_302 = 4'h1 == _T_1277 ? $signed(_T_1473_1) : $signed(_T_1473_0);
  assign _GEN_303 = 4'h2 == _T_1277 ? $signed(_T_1473_2) : $signed(_GEN_302);
  assign _GEN_304 = 4'h3 == _T_1277 ? $signed(_T_1473_3) : $signed(_GEN_303);
  assign _GEN_305 = 4'h4 == _T_1277 ? $signed(_T_1473_4) : $signed(_GEN_304);
  assign _GEN_306 = 4'h5 == _T_1277 ? $signed(_T_1473_5) : $signed(_GEN_305);
  assign _GEN_307 = 4'h6 == _T_1277 ? $signed(_T_1473_6) : $signed(_GEN_306);
  assign _GEN_308 = 4'h7 == _T_1277 ? $signed(_T_1473_7) : $signed(_GEN_307);
  assign _GEN_309 = 4'h8 == _T_1277 ? $signed(_T_1473_8) : $signed(_GEN_308);
  assign _GEN_310 = 4'h9 == _T_1277 ? $signed(_T_1473_9) : $signed(_GEN_309);
  assign _GEN_311 = 4'ha == _T_1277 ? $signed(_T_1473_10) : $signed(_GEN_310);
  assign _GEN_312 = 4'hb == _T_1277 ? $signed(_T_1473_11) : $signed(_GEN_311);
  assign _GEN_313 = 4'hc == _T_1277 ? $signed(_T_1473_12) : $signed(_GEN_312);
  assign _GEN_314 = 4'hd == _T_1277 ? $signed(_T_1473_13) : $signed(_GEN_313);
  assign _GEN_315 = 4'he == _T_1277 ? $signed(_T_1473_14) : $signed(_GEN_314);
  assign _GEN_316 = 4'hf == _T_1277 ? $signed(_T_1473_15) : $signed(_GEN_315);
  assign _GEN_19 = _GEN_331;
  assign _GEN_317 = 4'h1 == _T_1278 ? $signed(_T_1543_1) : $signed(_T_1543_0);
  assign _GEN_318 = 4'h2 == _T_1278 ? $signed(_T_1543_2) : $signed(_GEN_317);
  assign _GEN_319 = 4'h3 == _T_1278 ? $signed(_T_1543_3) : $signed(_GEN_318);
  assign _GEN_320 = 4'h4 == _T_1278 ? $signed(_T_1543_4) : $signed(_GEN_319);
  assign _GEN_321 = 4'h5 == _T_1278 ? $signed(_T_1543_5) : $signed(_GEN_320);
  assign _GEN_322 = 4'h6 == _T_1278 ? $signed(_T_1543_6) : $signed(_GEN_321);
  assign _GEN_323 = 4'h7 == _T_1278 ? $signed(_T_1543_7) : $signed(_GEN_322);
  assign _GEN_324 = 4'h8 == _T_1278 ? $signed(_T_1543_8) : $signed(_GEN_323);
  assign _GEN_325 = 4'h9 == _T_1278 ? $signed(_T_1543_9) : $signed(_GEN_324);
  assign _GEN_326 = 4'ha == _T_1278 ? $signed(_T_1543_10) : $signed(_GEN_325);
  assign _GEN_327 = 4'hb == _T_1278 ? $signed(_T_1543_11) : $signed(_GEN_326);
  assign _GEN_328 = 4'hc == _T_1278 ? $signed(_T_1543_12) : $signed(_GEN_327);
  assign _GEN_329 = 4'hd == _T_1278 ? $signed(_T_1543_13) : $signed(_GEN_328);
  assign _GEN_330 = 4'he == _T_1278 ? $signed(_T_1543_14) : $signed(_GEN_329);
  assign _GEN_331 = 4'hf == _T_1278 ? $signed(_T_1543_15) : $signed(_GEN_330);
  assign _T_1846 = $signed(_GEN_18) + $signed(_GEN_19);
  assign _T_1847 = _T_1846[5:0];
  assign _T_1848 = $signed(_T_1847);
  assign _GEN_20 = _GEN_346;
  assign _GEN_332 = 4'h1 == _T_1279 ? $signed(_T_1613_1) : $signed(_T_1613_0);
  assign _GEN_333 = 4'h2 == _T_1279 ? $signed(_T_1613_2) : $signed(_GEN_332);
  assign _GEN_334 = 4'h3 == _T_1279 ? $signed(_T_1613_3) : $signed(_GEN_333);
  assign _GEN_335 = 4'h4 == _T_1279 ? $signed(_T_1613_4) : $signed(_GEN_334);
  assign _GEN_336 = 4'h5 == _T_1279 ? $signed(_T_1613_5) : $signed(_GEN_335);
  assign _GEN_337 = 4'h6 == _T_1279 ? $signed(_T_1613_6) : $signed(_GEN_336);
  assign _GEN_338 = 4'h7 == _T_1279 ? $signed(_T_1613_7) : $signed(_GEN_337);
  assign _GEN_339 = 4'h8 == _T_1279 ? $signed(_T_1613_8) : $signed(_GEN_338);
  assign _GEN_340 = 4'h9 == _T_1279 ? $signed(_T_1613_9) : $signed(_GEN_339);
  assign _GEN_341 = 4'ha == _T_1279 ? $signed(_T_1613_10) : $signed(_GEN_340);
  assign _GEN_342 = 4'hb == _T_1279 ? $signed(_T_1613_11) : $signed(_GEN_341);
  assign _GEN_343 = 4'hc == _T_1279 ? $signed(_T_1613_12) : $signed(_GEN_342);
  assign _GEN_344 = 4'hd == _T_1279 ? $signed(_T_1613_13) : $signed(_GEN_343);
  assign _GEN_345 = 4'he == _T_1279 ? $signed(_T_1613_14) : $signed(_GEN_344);
  assign _GEN_346 = 4'hf == _T_1279 ? $signed(_T_1613_15) : $signed(_GEN_345);
  assign _GEN_21 = _GEN_361;
  assign _GEN_347 = 4'h1 == _T_1280 ? $signed(_T_1683_1) : $signed(_T_1683_0);
  assign _GEN_348 = 4'h2 == _T_1280 ? $signed(_T_1683_2) : $signed(_GEN_347);
  assign _GEN_349 = 4'h3 == _T_1280 ? $signed(_T_1683_3) : $signed(_GEN_348);
  assign _GEN_350 = 4'h4 == _T_1280 ? $signed(_T_1683_4) : $signed(_GEN_349);
  assign _GEN_351 = 4'h5 == _T_1280 ? $signed(_T_1683_5) : $signed(_GEN_350);
  assign _GEN_352 = 4'h6 == _T_1280 ? $signed(_T_1683_6) : $signed(_GEN_351);
  assign _GEN_353 = 4'h7 == _T_1280 ? $signed(_T_1683_7) : $signed(_GEN_352);
  assign _GEN_354 = 4'h8 == _T_1280 ? $signed(_T_1683_8) : $signed(_GEN_353);
  assign _GEN_355 = 4'h9 == _T_1280 ? $signed(_T_1683_9) : $signed(_GEN_354);
  assign _GEN_356 = 4'ha == _T_1280 ? $signed(_T_1683_10) : $signed(_GEN_355);
  assign _GEN_357 = 4'hb == _T_1280 ? $signed(_T_1683_11) : $signed(_GEN_356);
  assign _GEN_358 = 4'hc == _T_1280 ? $signed(_T_1683_12) : $signed(_GEN_357);
  assign _GEN_359 = 4'hd == _T_1280 ? $signed(_T_1683_13) : $signed(_GEN_358);
  assign _GEN_360 = 4'he == _T_1280 ? $signed(_T_1683_14) : $signed(_GEN_359);
  assign _GEN_361 = 4'hf == _T_1280 ? $signed(_T_1683_15) : $signed(_GEN_360);
  assign _T_1849 = $signed(_GEN_20) + $signed(_GEN_21);
  assign _T_1850 = _T_1849[5:0];
  assign _T_1851 = $signed(_T_1850);
  assign _GEN_22 = _GEN_376;
  assign _GEN_362 = 4'h1 == _T_1281 ? $signed(_T_1753_1) : $signed(_T_1753_0);
  assign _GEN_363 = 4'h2 == _T_1281 ? $signed(_T_1753_2) : $signed(_GEN_362);
  assign _GEN_364 = 4'h3 == _T_1281 ? $signed(_T_1753_3) : $signed(_GEN_363);
  assign _GEN_365 = 4'h4 == _T_1281 ? $signed(_T_1753_4) : $signed(_GEN_364);
  assign _GEN_366 = 4'h5 == _T_1281 ? $signed(_T_1753_5) : $signed(_GEN_365);
  assign _GEN_367 = 4'h6 == _T_1281 ? $signed(_T_1753_6) : $signed(_GEN_366);
  assign _GEN_368 = 4'h7 == _T_1281 ? $signed(_T_1753_7) : $signed(_GEN_367);
  assign _GEN_369 = 4'h8 == _T_1281 ? $signed(_T_1753_8) : $signed(_GEN_368);
  assign _GEN_370 = 4'h9 == _T_1281 ? $signed(_T_1753_9) : $signed(_GEN_369);
  assign _GEN_371 = 4'ha == _T_1281 ? $signed(_T_1753_10) : $signed(_GEN_370);
  assign _GEN_372 = 4'hb == _T_1281 ? $signed(_T_1753_11) : $signed(_GEN_371);
  assign _GEN_373 = 4'hc == _T_1281 ? $signed(_T_1753_12) : $signed(_GEN_372);
  assign _GEN_374 = 4'hd == _T_1281 ? $signed(_T_1753_13) : $signed(_GEN_373);
  assign _GEN_375 = 4'he == _T_1281 ? $signed(_T_1753_14) : $signed(_GEN_374);
  assign _GEN_376 = 4'hf == _T_1281 ? $signed(_T_1753_15) : $signed(_GEN_375);
  assign _GEN_23 = _GEN_391;
  assign _GEN_377 = 4'h1 == _T_1282 ? $signed(_T_1823_1) : $signed(_T_1823_0);
  assign _GEN_378 = 4'h2 == _T_1282 ? $signed(_T_1823_2) : $signed(_GEN_377);
  assign _GEN_379 = 4'h3 == _T_1282 ? $signed(_T_1823_3) : $signed(_GEN_378);
  assign _GEN_380 = 4'h4 == _T_1282 ? $signed(_T_1823_4) : $signed(_GEN_379);
  assign _GEN_381 = 4'h5 == _T_1282 ? $signed(_T_1823_5) : $signed(_GEN_380);
  assign _GEN_382 = 4'h6 == _T_1282 ? $signed(_T_1823_6) : $signed(_GEN_381);
  assign _GEN_383 = 4'h7 == _T_1282 ? $signed(_T_1823_7) : $signed(_GEN_382);
  assign _GEN_384 = 4'h8 == _T_1282 ? $signed(_T_1823_8) : $signed(_GEN_383);
  assign _GEN_385 = 4'h9 == _T_1282 ? $signed(_T_1823_9) : $signed(_GEN_384);
  assign _GEN_386 = 4'ha == _T_1282 ? $signed(_T_1823_10) : $signed(_GEN_385);
  assign _GEN_387 = 4'hb == _T_1282 ? $signed(_T_1823_11) : $signed(_GEN_386);
  assign _GEN_388 = 4'hc == _T_1282 ? $signed(_T_1823_12) : $signed(_GEN_387);
  assign _GEN_389 = 4'hd == _T_1282 ? $signed(_T_1823_13) : $signed(_GEN_388);
  assign _GEN_390 = 4'he == _T_1282 ? $signed(_T_1823_14) : $signed(_GEN_389);
  assign _GEN_391 = 4'hf == _T_1282 ? $signed(_T_1823_15) : $signed(_GEN_390);
  assign _T_1852 = $signed(_GEN_22) + $signed(_GEN_23);
  assign _T_1853 = _T_1852[5:0];
  assign _T_1854 = $signed(_T_1853);
  assign _T_1855 = $signed(_T_1845) + $signed(_T_1848);
  assign _T_1856 = _T_1855[5:0];
  assign _T_1857 = $signed(_T_1856);
  assign _T_1858 = $signed(_T_1851) + $signed(_T_1854);
  assign _T_1859 = _T_1858[5:0];
  assign _T_1860 = $signed(_T_1859);
  assign _T_1861 = $signed(_T_1857) + $signed(_T_1860);
  assign _T_1862 = _T_1861[5:0];
  assign _T_1863 = $signed(_T_1862);
  assign MulAdd_2_io_a = _T_1868;
  assign MulAdd_2_io_b = $signed(_GEN_514);
  assign MulAdd_2_io_m = mean_io_output;
  assign MulAdd_2_io_c = _T_1870;
  assign _T_1865 = mem_io_out[63:32];
  assign _T_1866 = io_memSel ? 32'h0 : _T_1865;
  assign _T_1867 = _T_1866[31:16];
  assign _T_1868 = $signed(_T_1867);
  assign _T_1869 = _T_1866[15:0];
  assign _T_1870 = $signed(_T_1869);
  assign signs_2 = MulAdd_2_io_r[31];
  assign Accumulator_3_clock = clock;
  assign Accumulator_3_io_in = {{26{_T_2459[5]}},_T_2459};
  assign Accumulator_3_io_sel = io_accSel;
  assign Accumulator_3_io_en = io_accEn;
  assign Accumulator_3_io_reset = io_accReset;
  assign _T_1871 = xnor$_io_out_3[3:0];
  assign _T_1872 = xnor$_io_out_3[7:4];
  assign _T_1873 = xnor$_io_out_3[11:8];
  assign _T_1874 = xnor$_io_out_3[15:12];
  assign _T_1875 = xnor$_io_out_3[19:16];
  assign _T_1876 = xnor$_io_out_3[23:20];
  assign _T_1877 = xnor$_io_out_3[27:24];
  assign _T_1878 = xnor$_io_out_3[31:28];
  assign _T_1929_0 = _T_1881;
  assign _T_1929_1 = _T_1884;
  assign _T_1929_2 = _T_1887;
  assign _T_1929_3 = _T_1890;
  assign _T_1929_4 = _T_1893;
  assign _T_1929_5 = _T_1896;
  assign _T_1929_6 = _T_1899;
  assign _T_1929_7 = _T_1902;
  assign _T_1929_8 = _T_1905;
  assign _T_1929_9 = _T_1908;
  assign _T_1929_10 = _T_1911;
  assign _T_1929_11 = _T_1914;
  assign _T_1929_12 = _T_1917;
  assign _T_1929_13 = _T_1920;
  assign _T_1929_14 = _T_1923;
  assign _T_1929_15 = _T_1926;
  assign _T_1999_0 = _T_1951;
  assign _T_1999_1 = _T_1954;
  assign _T_1999_2 = _T_1957;
  assign _T_1999_3 = _T_1960;
  assign _T_1999_4 = _T_1963;
  assign _T_1999_5 = _T_1966;
  assign _T_1999_6 = _T_1969;
  assign _T_1999_7 = _T_1972;
  assign _T_1999_8 = _T_1975;
  assign _T_1999_9 = _T_1978;
  assign _T_1999_10 = _T_1981;
  assign _T_1999_11 = _T_1984;
  assign _T_1999_12 = _T_1987;
  assign _T_1999_13 = _T_1990;
  assign _T_1999_14 = _T_1993;
  assign _T_1999_15 = _T_1996;
  assign _T_2069_0 = _T_2021;
  assign _T_2069_1 = _T_2024;
  assign _T_2069_2 = _T_2027;
  assign _T_2069_3 = _T_2030;
  assign _T_2069_4 = _T_2033;
  assign _T_2069_5 = _T_2036;
  assign _T_2069_6 = _T_2039;
  assign _T_2069_7 = _T_2042;
  assign _T_2069_8 = _T_2045;
  assign _T_2069_9 = _T_2048;
  assign _T_2069_10 = _T_2051;
  assign _T_2069_11 = _T_2054;
  assign _T_2069_12 = _T_2057;
  assign _T_2069_13 = _T_2060;
  assign _T_2069_14 = _T_2063;
  assign _T_2069_15 = _T_2066;
  assign _T_2139_0 = _T_2091;
  assign _T_2139_1 = _T_2094;
  assign _T_2139_2 = _T_2097;
  assign _T_2139_3 = _T_2100;
  assign _T_2139_4 = _T_2103;
  assign _T_2139_5 = _T_2106;
  assign _T_2139_6 = _T_2109;
  assign _T_2139_7 = _T_2112;
  assign _T_2139_8 = _T_2115;
  assign _T_2139_9 = _T_2118;
  assign _T_2139_10 = _T_2121;
  assign _T_2139_11 = _T_2124;
  assign _T_2139_12 = _T_2127;
  assign _T_2139_13 = _T_2130;
  assign _T_2139_14 = _T_2133;
  assign _T_2139_15 = _T_2136;
  assign _T_2209_0 = _T_2161;
  assign _T_2209_1 = _T_2164;
  assign _T_2209_2 = _T_2167;
  assign _T_2209_3 = _T_2170;
  assign _T_2209_4 = _T_2173;
  assign _T_2209_5 = _T_2176;
  assign _T_2209_6 = _T_2179;
  assign _T_2209_7 = _T_2182;
  assign _T_2209_8 = _T_2185;
  assign _T_2209_9 = _T_2188;
  assign _T_2209_10 = _T_2191;
  assign _T_2209_11 = _T_2194;
  assign _T_2209_12 = _T_2197;
  assign _T_2209_13 = _T_2200;
  assign _T_2209_14 = _T_2203;
  assign _T_2209_15 = _T_2206;
  assign _T_2279_0 = _T_2231;
  assign _T_2279_1 = _T_2234;
  assign _T_2279_2 = _T_2237;
  assign _T_2279_3 = _T_2240;
  assign _T_2279_4 = _T_2243;
  assign _T_2279_5 = _T_2246;
  assign _T_2279_6 = _T_2249;
  assign _T_2279_7 = _T_2252;
  assign _T_2279_8 = _T_2255;
  assign _T_2279_9 = _T_2258;
  assign _T_2279_10 = _T_2261;
  assign _T_2279_11 = _T_2264;
  assign _T_2279_12 = _T_2267;
  assign _T_2279_13 = _T_2270;
  assign _T_2279_14 = _T_2273;
  assign _T_2279_15 = _T_2276;
  assign _T_2349_0 = _T_2301;
  assign _T_2349_1 = _T_2304;
  assign _T_2349_2 = _T_2307;
  assign _T_2349_3 = _T_2310;
  assign _T_2349_4 = _T_2313;
  assign _T_2349_5 = _T_2316;
  assign _T_2349_6 = _T_2319;
  assign _T_2349_7 = _T_2322;
  assign _T_2349_8 = _T_2325;
  assign _T_2349_9 = _T_2328;
  assign _T_2349_10 = _T_2331;
  assign _T_2349_11 = _T_2334;
  assign _T_2349_12 = _T_2337;
  assign _T_2349_13 = _T_2340;
  assign _T_2349_14 = _T_2343;
  assign _T_2349_15 = _T_2346;
  assign _T_2419_0 = _T_2371;
  assign _T_2419_1 = _T_2374;
  assign _T_2419_2 = _T_2377;
  assign _T_2419_3 = _T_2380;
  assign _T_2419_4 = _T_2383;
  assign _T_2419_5 = _T_2386;
  assign _T_2419_6 = _T_2389;
  assign _T_2419_7 = _T_2392;
  assign _T_2419_8 = _T_2395;
  assign _T_2419_9 = _T_2398;
  assign _T_2419_10 = _T_2401;
  assign _T_2419_11 = _T_2404;
  assign _T_2419_12 = _T_2407;
  assign _T_2419_13 = _T_2410;
  assign _T_2419_14 = _T_2413;
  assign _T_2419_15 = _T_2416;
  assign _GEN_24 = _GEN_406;
  assign _GEN_392 = 4'h1 == _T_1871 ? $signed(_T_1929_1) : $signed(_T_1929_0);
  assign _GEN_393 = 4'h2 == _T_1871 ? $signed(_T_1929_2) : $signed(_GEN_392);
  assign _GEN_394 = 4'h3 == _T_1871 ? $signed(_T_1929_3) : $signed(_GEN_393);
  assign _GEN_395 = 4'h4 == _T_1871 ? $signed(_T_1929_4) : $signed(_GEN_394);
  assign _GEN_396 = 4'h5 == _T_1871 ? $signed(_T_1929_5) : $signed(_GEN_395);
  assign _GEN_397 = 4'h6 == _T_1871 ? $signed(_T_1929_6) : $signed(_GEN_396);
  assign _GEN_398 = 4'h7 == _T_1871 ? $signed(_T_1929_7) : $signed(_GEN_397);
  assign _GEN_399 = 4'h8 == _T_1871 ? $signed(_T_1929_8) : $signed(_GEN_398);
  assign _GEN_400 = 4'h9 == _T_1871 ? $signed(_T_1929_9) : $signed(_GEN_399);
  assign _GEN_401 = 4'ha == _T_1871 ? $signed(_T_1929_10) : $signed(_GEN_400);
  assign _GEN_402 = 4'hb == _T_1871 ? $signed(_T_1929_11) : $signed(_GEN_401);
  assign _GEN_403 = 4'hc == _T_1871 ? $signed(_T_1929_12) : $signed(_GEN_402);
  assign _GEN_404 = 4'hd == _T_1871 ? $signed(_T_1929_13) : $signed(_GEN_403);
  assign _GEN_405 = 4'he == _T_1871 ? $signed(_T_1929_14) : $signed(_GEN_404);
  assign _GEN_406 = 4'hf == _T_1871 ? $signed(_T_1929_15) : $signed(_GEN_405);
  assign _GEN_25 = _GEN_421;
  assign _GEN_407 = 4'h1 == _T_1872 ? $signed(_T_1999_1) : $signed(_T_1999_0);
  assign _GEN_408 = 4'h2 == _T_1872 ? $signed(_T_1999_2) : $signed(_GEN_407);
  assign _GEN_409 = 4'h3 == _T_1872 ? $signed(_T_1999_3) : $signed(_GEN_408);
  assign _GEN_410 = 4'h4 == _T_1872 ? $signed(_T_1999_4) : $signed(_GEN_409);
  assign _GEN_411 = 4'h5 == _T_1872 ? $signed(_T_1999_5) : $signed(_GEN_410);
  assign _GEN_412 = 4'h6 == _T_1872 ? $signed(_T_1999_6) : $signed(_GEN_411);
  assign _GEN_413 = 4'h7 == _T_1872 ? $signed(_T_1999_7) : $signed(_GEN_412);
  assign _GEN_414 = 4'h8 == _T_1872 ? $signed(_T_1999_8) : $signed(_GEN_413);
  assign _GEN_415 = 4'h9 == _T_1872 ? $signed(_T_1999_9) : $signed(_GEN_414);
  assign _GEN_416 = 4'ha == _T_1872 ? $signed(_T_1999_10) : $signed(_GEN_415);
  assign _GEN_417 = 4'hb == _T_1872 ? $signed(_T_1999_11) : $signed(_GEN_416);
  assign _GEN_418 = 4'hc == _T_1872 ? $signed(_T_1999_12) : $signed(_GEN_417);
  assign _GEN_419 = 4'hd == _T_1872 ? $signed(_T_1999_13) : $signed(_GEN_418);
  assign _GEN_420 = 4'he == _T_1872 ? $signed(_T_1999_14) : $signed(_GEN_419);
  assign _GEN_421 = 4'hf == _T_1872 ? $signed(_T_1999_15) : $signed(_GEN_420);
  assign _T_2439 = $signed(_GEN_24) + $signed(_GEN_25);
  assign _T_2440 = _T_2439[5:0];
  assign _T_2441 = $signed(_T_2440);
  assign _GEN_26 = _GEN_436;
  assign _GEN_422 = 4'h1 == _T_1873 ? $signed(_T_2069_1) : $signed(_T_2069_0);
  assign _GEN_423 = 4'h2 == _T_1873 ? $signed(_T_2069_2) : $signed(_GEN_422);
  assign _GEN_424 = 4'h3 == _T_1873 ? $signed(_T_2069_3) : $signed(_GEN_423);
  assign _GEN_425 = 4'h4 == _T_1873 ? $signed(_T_2069_4) : $signed(_GEN_424);
  assign _GEN_426 = 4'h5 == _T_1873 ? $signed(_T_2069_5) : $signed(_GEN_425);
  assign _GEN_427 = 4'h6 == _T_1873 ? $signed(_T_2069_6) : $signed(_GEN_426);
  assign _GEN_428 = 4'h7 == _T_1873 ? $signed(_T_2069_7) : $signed(_GEN_427);
  assign _GEN_429 = 4'h8 == _T_1873 ? $signed(_T_2069_8) : $signed(_GEN_428);
  assign _GEN_430 = 4'h9 == _T_1873 ? $signed(_T_2069_9) : $signed(_GEN_429);
  assign _GEN_431 = 4'ha == _T_1873 ? $signed(_T_2069_10) : $signed(_GEN_430);
  assign _GEN_432 = 4'hb == _T_1873 ? $signed(_T_2069_11) : $signed(_GEN_431);
  assign _GEN_433 = 4'hc == _T_1873 ? $signed(_T_2069_12) : $signed(_GEN_432);
  assign _GEN_434 = 4'hd == _T_1873 ? $signed(_T_2069_13) : $signed(_GEN_433);
  assign _GEN_435 = 4'he == _T_1873 ? $signed(_T_2069_14) : $signed(_GEN_434);
  assign _GEN_436 = 4'hf == _T_1873 ? $signed(_T_2069_15) : $signed(_GEN_435);
  assign _GEN_27 = _GEN_451;
  assign _GEN_437 = 4'h1 == _T_1874 ? $signed(_T_2139_1) : $signed(_T_2139_0);
  assign _GEN_438 = 4'h2 == _T_1874 ? $signed(_T_2139_2) : $signed(_GEN_437);
  assign _GEN_439 = 4'h3 == _T_1874 ? $signed(_T_2139_3) : $signed(_GEN_438);
  assign _GEN_440 = 4'h4 == _T_1874 ? $signed(_T_2139_4) : $signed(_GEN_439);
  assign _GEN_441 = 4'h5 == _T_1874 ? $signed(_T_2139_5) : $signed(_GEN_440);
  assign _GEN_442 = 4'h6 == _T_1874 ? $signed(_T_2139_6) : $signed(_GEN_441);
  assign _GEN_443 = 4'h7 == _T_1874 ? $signed(_T_2139_7) : $signed(_GEN_442);
  assign _GEN_444 = 4'h8 == _T_1874 ? $signed(_T_2139_8) : $signed(_GEN_443);
  assign _GEN_445 = 4'h9 == _T_1874 ? $signed(_T_2139_9) : $signed(_GEN_444);
  assign _GEN_446 = 4'ha == _T_1874 ? $signed(_T_2139_10) : $signed(_GEN_445);
  assign _GEN_447 = 4'hb == _T_1874 ? $signed(_T_2139_11) : $signed(_GEN_446);
  assign _GEN_448 = 4'hc == _T_1874 ? $signed(_T_2139_12) : $signed(_GEN_447);
  assign _GEN_449 = 4'hd == _T_1874 ? $signed(_T_2139_13) : $signed(_GEN_448);
  assign _GEN_450 = 4'he == _T_1874 ? $signed(_T_2139_14) : $signed(_GEN_449);
  assign _GEN_451 = 4'hf == _T_1874 ? $signed(_T_2139_15) : $signed(_GEN_450);
  assign _T_2442 = $signed(_GEN_26) + $signed(_GEN_27);
  assign _T_2443 = _T_2442[5:0];
  assign _T_2444 = $signed(_T_2443);
  assign _GEN_28 = _GEN_466;
  assign _GEN_452 = 4'h1 == _T_1875 ? $signed(_T_2209_1) : $signed(_T_2209_0);
  assign _GEN_453 = 4'h2 == _T_1875 ? $signed(_T_2209_2) : $signed(_GEN_452);
  assign _GEN_454 = 4'h3 == _T_1875 ? $signed(_T_2209_3) : $signed(_GEN_453);
  assign _GEN_455 = 4'h4 == _T_1875 ? $signed(_T_2209_4) : $signed(_GEN_454);
  assign _GEN_456 = 4'h5 == _T_1875 ? $signed(_T_2209_5) : $signed(_GEN_455);
  assign _GEN_457 = 4'h6 == _T_1875 ? $signed(_T_2209_6) : $signed(_GEN_456);
  assign _GEN_458 = 4'h7 == _T_1875 ? $signed(_T_2209_7) : $signed(_GEN_457);
  assign _GEN_459 = 4'h8 == _T_1875 ? $signed(_T_2209_8) : $signed(_GEN_458);
  assign _GEN_460 = 4'h9 == _T_1875 ? $signed(_T_2209_9) : $signed(_GEN_459);
  assign _GEN_461 = 4'ha == _T_1875 ? $signed(_T_2209_10) : $signed(_GEN_460);
  assign _GEN_462 = 4'hb == _T_1875 ? $signed(_T_2209_11) : $signed(_GEN_461);
  assign _GEN_463 = 4'hc == _T_1875 ? $signed(_T_2209_12) : $signed(_GEN_462);
  assign _GEN_464 = 4'hd == _T_1875 ? $signed(_T_2209_13) : $signed(_GEN_463);
  assign _GEN_465 = 4'he == _T_1875 ? $signed(_T_2209_14) : $signed(_GEN_464);
  assign _GEN_466 = 4'hf == _T_1875 ? $signed(_T_2209_15) : $signed(_GEN_465);
  assign _GEN_29 = _GEN_481;
  assign _GEN_467 = 4'h1 == _T_1876 ? $signed(_T_2279_1) : $signed(_T_2279_0);
  assign _GEN_468 = 4'h2 == _T_1876 ? $signed(_T_2279_2) : $signed(_GEN_467);
  assign _GEN_469 = 4'h3 == _T_1876 ? $signed(_T_2279_3) : $signed(_GEN_468);
  assign _GEN_470 = 4'h4 == _T_1876 ? $signed(_T_2279_4) : $signed(_GEN_469);
  assign _GEN_471 = 4'h5 == _T_1876 ? $signed(_T_2279_5) : $signed(_GEN_470);
  assign _GEN_472 = 4'h6 == _T_1876 ? $signed(_T_2279_6) : $signed(_GEN_471);
  assign _GEN_473 = 4'h7 == _T_1876 ? $signed(_T_2279_7) : $signed(_GEN_472);
  assign _GEN_474 = 4'h8 == _T_1876 ? $signed(_T_2279_8) : $signed(_GEN_473);
  assign _GEN_475 = 4'h9 == _T_1876 ? $signed(_T_2279_9) : $signed(_GEN_474);
  assign _GEN_476 = 4'ha == _T_1876 ? $signed(_T_2279_10) : $signed(_GEN_475);
  assign _GEN_477 = 4'hb == _T_1876 ? $signed(_T_2279_11) : $signed(_GEN_476);
  assign _GEN_478 = 4'hc == _T_1876 ? $signed(_T_2279_12) : $signed(_GEN_477);
  assign _GEN_479 = 4'hd == _T_1876 ? $signed(_T_2279_13) : $signed(_GEN_478);
  assign _GEN_480 = 4'he == _T_1876 ? $signed(_T_2279_14) : $signed(_GEN_479);
  assign _GEN_481 = 4'hf == _T_1876 ? $signed(_T_2279_15) : $signed(_GEN_480);
  assign _T_2445 = $signed(_GEN_28) + $signed(_GEN_29);
  assign _T_2446 = _T_2445[5:0];
  assign _T_2447 = $signed(_T_2446);
  assign _GEN_30 = _GEN_496;
  assign _GEN_482 = 4'h1 == _T_1877 ? $signed(_T_2349_1) : $signed(_T_2349_0);
  assign _GEN_483 = 4'h2 == _T_1877 ? $signed(_T_2349_2) : $signed(_GEN_482);
  assign _GEN_484 = 4'h3 == _T_1877 ? $signed(_T_2349_3) : $signed(_GEN_483);
  assign _GEN_485 = 4'h4 == _T_1877 ? $signed(_T_2349_4) : $signed(_GEN_484);
  assign _GEN_486 = 4'h5 == _T_1877 ? $signed(_T_2349_5) : $signed(_GEN_485);
  assign _GEN_487 = 4'h6 == _T_1877 ? $signed(_T_2349_6) : $signed(_GEN_486);
  assign _GEN_488 = 4'h7 == _T_1877 ? $signed(_T_2349_7) : $signed(_GEN_487);
  assign _GEN_489 = 4'h8 == _T_1877 ? $signed(_T_2349_8) : $signed(_GEN_488);
  assign _GEN_490 = 4'h9 == _T_1877 ? $signed(_T_2349_9) : $signed(_GEN_489);
  assign _GEN_491 = 4'ha == _T_1877 ? $signed(_T_2349_10) : $signed(_GEN_490);
  assign _GEN_492 = 4'hb == _T_1877 ? $signed(_T_2349_11) : $signed(_GEN_491);
  assign _GEN_493 = 4'hc == _T_1877 ? $signed(_T_2349_12) : $signed(_GEN_492);
  assign _GEN_494 = 4'hd == _T_1877 ? $signed(_T_2349_13) : $signed(_GEN_493);
  assign _GEN_495 = 4'he == _T_1877 ? $signed(_T_2349_14) : $signed(_GEN_494);
  assign _GEN_496 = 4'hf == _T_1877 ? $signed(_T_2349_15) : $signed(_GEN_495);
  assign _GEN_31 = _GEN_511;
  assign _GEN_497 = 4'h1 == _T_1878 ? $signed(_T_2419_1) : $signed(_T_2419_0);
  assign _GEN_498 = 4'h2 == _T_1878 ? $signed(_T_2419_2) : $signed(_GEN_497);
  assign _GEN_499 = 4'h3 == _T_1878 ? $signed(_T_2419_3) : $signed(_GEN_498);
  assign _GEN_500 = 4'h4 == _T_1878 ? $signed(_T_2419_4) : $signed(_GEN_499);
  assign _GEN_501 = 4'h5 == _T_1878 ? $signed(_T_2419_5) : $signed(_GEN_500);
  assign _GEN_502 = 4'h6 == _T_1878 ? $signed(_T_2419_6) : $signed(_GEN_501);
  assign _GEN_503 = 4'h7 == _T_1878 ? $signed(_T_2419_7) : $signed(_GEN_502);
  assign _GEN_504 = 4'h8 == _T_1878 ? $signed(_T_2419_8) : $signed(_GEN_503);
  assign _GEN_505 = 4'h9 == _T_1878 ? $signed(_T_2419_9) : $signed(_GEN_504);
  assign _GEN_506 = 4'ha == _T_1878 ? $signed(_T_2419_10) : $signed(_GEN_505);
  assign _GEN_507 = 4'hb == _T_1878 ? $signed(_T_2419_11) : $signed(_GEN_506);
  assign _GEN_508 = 4'hc == _T_1878 ? $signed(_T_2419_12) : $signed(_GEN_507);
  assign _GEN_509 = 4'hd == _T_1878 ? $signed(_T_2419_13) : $signed(_GEN_508);
  assign _GEN_510 = 4'he == _T_1878 ? $signed(_T_2419_14) : $signed(_GEN_509);
  assign _GEN_511 = 4'hf == _T_1878 ? $signed(_T_2419_15) : $signed(_GEN_510);
  assign _T_2448 = $signed(_GEN_30) + $signed(_GEN_31);
  assign _T_2449 = _T_2448[5:0];
  assign _T_2450 = $signed(_T_2449);
  assign _T_2451 = $signed(_T_2441) + $signed(_T_2444);
  assign _T_2452 = _T_2451[5:0];
  assign _T_2453 = $signed(_T_2452);
  assign _T_2454 = $signed(_T_2447) + $signed(_T_2450);
  assign _T_2455 = _T_2454[5:0];
  assign _T_2456 = $signed(_T_2455);
  assign _T_2457 = $signed(_T_2453) + $signed(_T_2456);
  assign _T_2458 = _T_2457[5:0];
  assign _T_2459 = $signed(_T_2458);
  assign MulAdd_3_io_a = _T_2464;
  assign MulAdd_3_io_b = $signed(_GEN_515);
  assign MulAdd_3_io_m = mean_io_output;
  assign MulAdd_3_io_c = _T_2466;
  assign _T_2461 = mem_io_out[31:0];
  assign _T_2462 = io_memSel ? 32'h0 : _T_2461;
  assign _T_2463 = _T_2462[31:16];
  assign _T_2464 = $signed(_T_2463);
  assign _T_2465 = _T_2462[15:0];
  assign _T_2466 = $signed(_T_2465);
  assign signs_3 = MulAdd_3_io_r[31];
  assign _T_2467 = {signs_2,signs_3};
  assign _T_2468 = {signs_0,signs_1};
  assign _T_2469 = {_T_2468,_T_2467};
  assign _GEN_512 = Accumulator_io_out[15:0];
  assign _GEN_513 = Accumulator_1_io_out[15:0];
  assign _GEN_514 = Accumulator_2_io_out[15:0];
  assign _GEN_515 = Accumulator_3_io_out[15:0];
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_516 = {1{$random}};
  _T_93 = _GEN_516[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_517 = {1{$random}};
  _T_96 = _GEN_517[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_518 = {1{$random}};
  _T_99 = _GEN_518[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_519 = {1{$random}};
  _T_102 = _GEN_519[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_520 = {1{$random}};
  _T_105 = _GEN_520[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_521 = {1{$random}};
  _T_108 = _GEN_521[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_522 = {1{$random}};
  _T_111 = _GEN_522[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_523 = {1{$random}};
  _T_114 = _GEN_523[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_524 = {1{$random}};
  _T_117 = _GEN_524[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_525 = {1{$random}};
  _T_120 = _GEN_525[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_526 = {1{$random}};
  _T_123 = _GEN_526[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_527 = {1{$random}};
  _T_126 = _GEN_527[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_528 = {1{$random}};
  _T_129 = _GEN_528[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_529 = {1{$random}};
  _T_132 = _GEN_529[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_530 = {1{$random}};
  _T_135 = _GEN_530[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_531 = {1{$random}};
  _T_138 = _GEN_531[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_532 = {1{$random}};
  _T_163 = _GEN_532[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_533 = {1{$random}};
  _T_166 = _GEN_533[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_534 = {1{$random}};
  _T_169 = _GEN_534[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_535 = {1{$random}};
  _T_172 = _GEN_535[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_536 = {1{$random}};
  _T_175 = _GEN_536[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_537 = {1{$random}};
  _T_178 = _GEN_537[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_538 = {1{$random}};
  _T_181 = _GEN_538[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_539 = {1{$random}};
  _T_184 = _GEN_539[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_540 = {1{$random}};
  _T_187 = _GEN_540[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_541 = {1{$random}};
  _T_190 = _GEN_541[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_542 = {1{$random}};
  _T_193 = _GEN_542[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_543 = {1{$random}};
  _T_196 = _GEN_543[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_544 = {1{$random}};
  _T_199 = _GEN_544[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_545 = {1{$random}};
  _T_202 = _GEN_545[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_546 = {1{$random}};
  _T_205 = _GEN_546[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_547 = {1{$random}};
  _T_208 = _GEN_547[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_548 = {1{$random}};
  _T_233 = _GEN_548[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_549 = {1{$random}};
  _T_236 = _GEN_549[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_550 = {1{$random}};
  _T_239 = _GEN_550[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_551 = {1{$random}};
  _T_242 = _GEN_551[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_552 = {1{$random}};
  _T_245 = _GEN_552[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_553 = {1{$random}};
  _T_248 = _GEN_553[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_554 = {1{$random}};
  _T_251 = _GEN_554[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_555 = {1{$random}};
  _T_254 = _GEN_555[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_556 = {1{$random}};
  _T_257 = _GEN_556[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_557 = {1{$random}};
  _T_260 = _GEN_557[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_558 = {1{$random}};
  _T_263 = _GEN_558[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_559 = {1{$random}};
  _T_266 = _GEN_559[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_560 = {1{$random}};
  _T_269 = _GEN_560[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_561 = {1{$random}};
  _T_272 = _GEN_561[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_562 = {1{$random}};
  _T_275 = _GEN_562[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_563 = {1{$random}};
  _T_278 = _GEN_563[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_564 = {1{$random}};
  _T_303 = _GEN_564[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_565 = {1{$random}};
  _T_306 = _GEN_565[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_566 = {1{$random}};
  _T_309 = _GEN_566[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_567 = {1{$random}};
  _T_312 = _GEN_567[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_568 = {1{$random}};
  _T_315 = _GEN_568[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_569 = {1{$random}};
  _T_318 = _GEN_569[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_570 = {1{$random}};
  _T_321 = _GEN_570[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_571 = {1{$random}};
  _T_324 = _GEN_571[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_572 = {1{$random}};
  _T_327 = _GEN_572[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_573 = {1{$random}};
  _T_330 = _GEN_573[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_574 = {1{$random}};
  _T_333 = _GEN_574[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_575 = {1{$random}};
  _T_336 = _GEN_575[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_576 = {1{$random}};
  _T_339 = _GEN_576[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_577 = {1{$random}};
  _T_342 = _GEN_577[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_578 = {1{$random}};
  _T_345 = _GEN_578[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_579 = {1{$random}};
  _T_348 = _GEN_579[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_580 = {1{$random}};
  _T_373 = _GEN_580[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_581 = {1{$random}};
  _T_376 = _GEN_581[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_582 = {1{$random}};
  _T_379 = _GEN_582[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_583 = {1{$random}};
  _T_382 = _GEN_583[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_584 = {1{$random}};
  _T_385 = _GEN_584[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_585 = {1{$random}};
  _T_388 = _GEN_585[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_586 = {1{$random}};
  _T_391 = _GEN_586[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_587 = {1{$random}};
  _T_394 = _GEN_587[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_588 = {1{$random}};
  _T_397 = _GEN_588[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_589 = {1{$random}};
  _T_400 = _GEN_589[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_590 = {1{$random}};
  _T_403 = _GEN_590[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_591 = {1{$random}};
  _T_406 = _GEN_591[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_592 = {1{$random}};
  _T_409 = _GEN_592[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_593 = {1{$random}};
  _T_412 = _GEN_593[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_594 = {1{$random}};
  _T_415 = _GEN_594[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_595 = {1{$random}};
  _T_418 = _GEN_595[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_596 = {1{$random}};
  _T_443 = _GEN_596[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_597 = {1{$random}};
  _T_446 = _GEN_597[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_598 = {1{$random}};
  _T_449 = _GEN_598[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_599 = {1{$random}};
  _T_452 = _GEN_599[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_600 = {1{$random}};
  _T_455 = _GEN_600[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_601 = {1{$random}};
  _T_458 = _GEN_601[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_602 = {1{$random}};
  _T_461 = _GEN_602[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_603 = {1{$random}};
  _T_464 = _GEN_603[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_604 = {1{$random}};
  _T_467 = _GEN_604[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_605 = {1{$random}};
  _T_470 = _GEN_605[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_606 = {1{$random}};
  _T_473 = _GEN_606[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_607 = {1{$random}};
  _T_476 = _GEN_607[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_608 = {1{$random}};
  _T_479 = _GEN_608[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_609 = {1{$random}};
  _T_482 = _GEN_609[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_610 = {1{$random}};
  _T_485 = _GEN_610[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_611 = {1{$random}};
  _T_488 = _GEN_611[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_612 = {1{$random}};
  _T_513 = _GEN_612[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_613 = {1{$random}};
  _T_516 = _GEN_613[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_614 = {1{$random}};
  _T_519 = _GEN_614[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_615 = {1{$random}};
  _T_522 = _GEN_615[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_616 = {1{$random}};
  _T_525 = _GEN_616[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_617 = {1{$random}};
  _T_528 = _GEN_617[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_618 = {1{$random}};
  _T_531 = _GEN_618[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_619 = {1{$random}};
  _T_534 = _GEN_619[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_620 = {1{$random}};
  _T_537 = _GEN_620[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_621 = {1{$random}};
  _T_540 = _GEN_621[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_622 = {1{$random}};
  _T_543 = _GEN_622[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_623 = {1{$random}};
  _T_546 = _GEN_623[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_624 = {1{$random}};
  _T_549 = _GEN_624[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_625 = {1{$random}};
  _T_552 = _GEN_625[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_626 = {1{$random}};
  _T_555 = _GEN_626[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_627 = {1{$random}};
  _T_558 = _GEN_627[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_628 = {1{$random}};
  _T_583 = _GEN_628[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_629 = {1{$random}};
  _T_586 = _GEN_629[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_630 = {1{$random}};
  _T_589 = _GEN_630[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_631 = {1{$random}};
  _T_592 = _GEN_631[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_632 = {1{$random}};
  _T_595 = _GEN_632[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_633 = {1{$random}};
  _T_598 = _GEN_633[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_634 = {1{$random}};
  _T_601 = _GEN_634[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_635 = {1{$random}};
  _T_604 = _GEN_635[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_636 = {1{$random}};
  _T_607 = _GEN_636[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_637 = {1{$random}};
  _T_610 = _GEN_637[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_638 = {1{$random}};
  _T_613 = _GEN_638[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_639 = {1{$random}};
  _T_616 = _GEN_639[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_640 = {1{$random}};
  _T_619 = _GEN_640[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_641 = {1{$random}};
  _T_622 = _GEN_641[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_642 = {1{$random}};
  _T_625 = _GEN_642[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_643 = {1{$random}};
  _T_628 = _GEN_643[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_644 = {1{$random}};
  _T_689 = _GEN_644[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_645 = {1{$random}};
  _T_692 = _GEN_645[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_646 = {1{$random}};
  _T_695 = _GEN_646[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_647 = {1{$random}};
  _T_698 = _GEN_647[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_648 = {1{$random}};
  _T_701 = _GEN_648[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_649 = {1{$random}};
  _T_704 = _GEN_649[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_650 = {1{$random}};
  _T_707 = _GEN_650[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_651 = {1{$random}};
  _T_710 = _GEN_651[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_652 = {1{$random}};
  _T_713 = _GEN_652[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_653 = {1{$random}};
  _T_716 = _GEN_653[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_654 = {1{$random}};
  _T_719 = _GEN_654[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_655 = {1{$random}};
  _T_722 = _GEN_655[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_656 = {1{$random}};
  _T_725 = _GEN_656[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_657 = {1{$random}};
  _T_728 = _GEN_657[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_658 = {1{$random}};
  _T_731 = _GEN_658[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_659 = {1{$random}};
  _T_734 = _GEN_659[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_660 = {1{$random}};
  _T_759 = _GEN_660[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_661 = {1{$random}};
  _T_762 = _GEN_661[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_662 = {1{$random}};
  _T_765 = _GEN_662[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_663 = {1{$random}};
  _T_768 = _GEN_663[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_664 = {1{$random}};
  _T_771 = _GEN_664[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_665 = {1{$random}};
  _T_774 = _GEN_665[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_666 = {1{$random}};
  _T_777 = _GEN_666[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_667 = {1{$random}};
  _T_780 = _GEN_667[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_668 = {1{$random}};
  _T_783 = _GEN_668[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_669 = {1{$random}};
  _T_786 = _GEN_669[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_670 = {1{$random}};
  _T_789 = _GEN_670[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_671 = {1{$random}};
  _T_792 = _GEN_671[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_672 = {1{$random}};
  _T_795 = _GEN_672[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_673 = {1{$random}};
  _T_798 = _GEN_673[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_674 = {1{$random}};
  _T_801 = _GEN_674[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_675 = {1{$random}};
  _T_804 = _GEN_675[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_676 = {1{$random}};
  _T_829 = _GEN_676[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_677 = {1{$random}};
  _T_832 = _GEN_677[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_678 = {1{$random}};
  _T_835 = _GEN_678[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_679 = {1{$random}};
  _T_838 = _GEN_679[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_680 = {1{$random}};
  _T_841 = _GEN_680[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_681 = {1{$random}};
  _T_844 = _GEN_681[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_682 = {1{$random}};
  _T_847 = _GEN_682[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_683 = {1{$random}};
  _T_850 = _GEN_683[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_684 = {1{$random}};
  _T_853 = _GEN_684[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_685 = {1{$random}};
  _T_856 = _GEN_685[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_686 = {1{$random}};
  _T_859 = _GEN_686[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_687 = {1{$random}};
  _T_862 = _GEN_687[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_688 = {1{$random}};
  _T_865 = _GEN_688[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_689 = {1{$random}};
  _T_868 = _GEN_689[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_690 = {1{$random}};
  _T_871 = _GEN_690[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_691 = {1{$random}};
  _T_874 = _GEN_691[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_692 = {1{$random}};
  _T_899 = _GEN_692[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_693 = {1{$random}};
  _T_902 = _GEN_693[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_694 = {1{$random}};
  _T_905 = _GEN_694[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_695 = {1{$random}};
  _T_908 = _GEN_695[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_696 = {1{$random}};
  _T_911 = _GEN_696[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_697 = {1{$random}};
  _T_914 = _GEN_697[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_698 = {1{$random}};
  _T_917 = _GEN_698[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_699 = {1{$random}};
  _T_920 = _GEN_699[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_700 = {1{$random}};
  _T_923 = _GEN_700[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_701 = {1{$random}};
  _T_926 = _GEN_701[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_702 = {1{$random}};
  _T_929 = _GEN_702[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_703 = {1{$random}};
  _T_932 = _GEN_703[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_704 = {1{$random}};
  _T_935 = _GEN_704[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_705 = {1{$random}};
  _T_938 = _GEN_705[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_706 = {1{$random}};
  _T_941 = _GEN_706[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_707 = {1{$random}};
  _T_944 = _GEN_707[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_708 = {1{$random}};
  _T_969 = _GEN_708[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_709 = {1{$random}};
  _T_972 = _GEN_709[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_710 = {1{$random}};
  _T_975 = _GEN_710[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_711 = {1{$random}};
  _T_978 = _GEN_711[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_712 = {1{$random}};
  _T_981 = _GEN_712[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_713 = {1{$random}};
  _T_984 = _GEN_713[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_714 = {1{$random}};
  _T_987 = _GEN_714[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_715 = {1{$random}};
  _T_990 = _GEN_715[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_716 = {1{$random}};
  _T_993 = _GEN_716[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_717 = {1{$random}};
  _T_996 = _GEN_717[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_718 = {1{$random}};
  _T_999 = _GEN_718[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_719 = {1{$random}};
  _T_1002 = _GEN_719[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_720 = {1{$random}};
  _T_1005 = _GEN_720[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_721 = {1{$random}};
  _T_1008 = _GEN_721[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_722 = {1{$random}};
  _T_1011 = _GEN_722[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_723 = {1{$random}};
  _T_1014 = _GEN_723[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_724 = {1{$random}};
  _T_1039 = _GEN_724[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_725 = {1{$random}};
  _T_1042 = _GEN_725[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_726 = {1{$random}};
  _T_1045 = _GEN_726[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_727 = {1{$random}};
  _T_1048 = _GEN_727[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_728 = {1{$random}};
  _T_1051 = _GEN_728[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_729 = {1{$random}};
  _T_1054 = _GEN_729[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_730 = {1{$random}};
  _T_1057 = _GEN_730[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_731 = {1{$random}};
  _T_1060 = _GEN_731[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_732 = {1{$random}};
  _T_1063 = _GEN_732[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_733 = {1{$random}};
  _T_1066 = _GEN_733[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_734 = {1{$random}};
  _T_1069 = _GEN_734[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_735 = {1{$random}};
  _T_1072 = _GEN_735[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_736 = {1{$random}};
  _T_1075 = _GEN_736[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_737 = {1{$random}};
  _T_1078 = _GEN_737[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_738 = {1{$random}};
  _T_1081 = _GEN_738[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_739 = {1{$random}};
  _T_1084 = _GEN_739[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_740 = {1{$random}};
  _T_1109 = _GEN_740[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_741 = {1{$random}};
  _T_1112 = _GEN_741[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_742 = {1{$random}};
  _T_1115 = _GEN_742[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_743 = {1{$random}};
  _T_1118 = _GEN_743[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_744 = {1{$random}};
  _T_1121 = _GEN_744[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_745 = {1{$random}};
  _T_1124 = _GEN_745[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_746 = {1{$random}};
  _T_1127 = _GEN_746[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_747 = {1{$random}};
  _T_1130 = _GEN_747[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_748 = {1{$random}};
  _T_1133 = _GEN_748[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_749 = {1{$random}};
  _T_1136 = _GEN_749[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_750 = {1{$random}};
  _T_1139 = _GEN_750[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_751 = {1{$random}};
  _T_1142 = _GEN_751[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_752 = {1{$random}};
  _T_1145 = _GEN_752[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_753 = {1{$random}};
  _T_1148 = _GEN_753[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_754 = {1{$random}};
  _T_1151 = _GEN_754[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_755 = {1{$random}};
  _T_1154 = _GEN_755[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_756 = {1{$random}};
  _T_1179 = _GEN_756[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_757 = {1{$random}};
  _T_1182 = _GEN_757[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_758 = {1{$random}};
  _T_1185 = _GEN_758[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_759 = {1{$random}};
  _T_1188 = _GEN_759[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_760 = {1{$random}};
  _T_1191 = _GEN_760[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_761 = {1{$random}};
  _T_1194 = _GEN_761[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_762 = {1{$random}};
  _T_1197 = _GEN_762[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_763 = {1{$random}};
  _T_1200 = _GEN_763[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_764 = {1{$random}};
  _T_1203 = _GEN_764[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_765 = {1{$random}};
  _T_1206 = _GEN_765[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_766 = {1{$random}};
  _T_1209 = _GEN_766[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_767 = {1{$random}};
  _T_1212 = _GEN_767[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_768 = {1{$random}};
  _T_1215 = _GEN_768[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_769 = {1{$random}};
  _T_1218 = _GEN_769[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_770 = {1{$random}};
  _T_1221 = _GEN_770[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_771 = {1{$random}};
  _T_1224 = _GEN_771[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_772 = {1{$random}};
  _T_1285 = _GEN_772[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_773 = {1{$random}};
  _T_1288 = _GEN_773[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_774 = {1{$random}};
  _T_1291 = _GEN_774[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_775 = {1{$random}};
  _T_1294 = _GEN_775[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_776 = {1{$random}};
  _T_1297 = _GEN_776[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_777 = {1{$random}};
  _T_1300 = _GEN_777[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_778 = {1{$random}};
  _T_1303 = _GEN_778[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_779 = {1{$random}};
  _T_1306 = _GEN_779[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_780 = {1{$random}};
  _T_1309 = _GEN_780[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_781 = {1{$random}};
  _T_1312 = _GEN_781[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_782 = {1{$random}};
  _T_1315 = _GEN_782[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_783 = {1{$random}};
  _T_1318 = _GEN_783[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_784 = {1{$random}};
  _T_1321 = _GEN_784[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_785 = {1{$random}};
  _T_1324 = _GEN_785[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_786 = {1{$random}};
  _T_1327 = _GEN_786[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_787 = {1{$random}};
  _T_1330 = _GEN_787[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_788 = {1{$random}};
  _T_1355 = _GEN_788[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_789 = {1{$random}};
  _T_1358 = _GEN_789[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_790 = {1{$random}};
  _T_1361 = _GEN_790[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_791 = {1{$random}};
  _T_1364 = _GEN_791[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_792 = {1{$random}};
  _T_1367 = _GEN_792[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_793 = {1{$random}};
  _T_1370 = _GEN_793[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_794 = {1{$random}};
  _T_1373 = _GEN_794[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_795 = {1{$random}};
  _T_1376 = _GEN_795[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_796 = {1{$random}};
  _T_1379 = _GEN_796[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_797 = {1{$random}};
  _T_1382 = _GEN_797[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_798 = {1{$random}};
  _T_1385 = _GEN_798[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_799 = {1{$random}};
  _T_1388 = _GEN_799[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_800 = {1{$random}};
  _T_1391 = _GEN_800[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_801 = {1{$random}};
  _T_1394 = _GEN_801[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_802 = {1{$random}};
  _T_1397 = _GEN_802[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_803 = {1{$random}};
  _T_1400 = _GEN_803[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_804 = {1{$random}};
  _T_1425 = _GEN_804[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_805 = {1{$random}};
  _T_1428 = _GEN_805[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_806 = {1{$random}};
  _T_1431 = _GEN_806[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_807 = {1{$random}};
  _T_1434 = _GEN_807[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_808 = {1{$random}};
  _T_1437 = _GEN_808[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_809 = {1{$random}};
  _T_1440 = _GEN_809[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_810 = {1{$random}};
  _T_1443 = _GEN_810[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_811 = {1{$random}};
  _T_1446 = _GEN_811[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_812 = {1{$random}};
  _T_1449 = _GEN_812[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_813 = {1{$random}};
  _T_1452 = _GEN_813[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_814 = {1{$random}};
  _T_1455 = _GEN_814[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_815 = {1{$random}};
  _T_1458 = _GEN_815[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_816 = {1{$random}};
  _T_1461 = _GEN_816[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_817 = {1{$random}};
  _T_1464 = _GEN_817[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_818 = {1{$random}};
  _T_1467 = _GEN_818[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_819 = {1{$random}};
  _T_1470 = _GEN_819[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_820 = {1{$random}};
  _T_1495 = _GEN_820[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_821 = {1{$random}};
  _T_1498 = _GEN_821[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_822 = {1{$random}};
  _T_1501 = _GEN_822[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_823 = {1{$random}};
  _T_1504 = _GEN_823[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_824 = {1{$random}};
  _T_1507 = _GEN_824[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_825 = {1{$random}};
  _T_1510 = _GEN_825[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_826 = {1{$random}};
  _T_1513 = _GEN_826[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_827 = {1{$random}};
  _T_1516 = _GEN_827[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_828 = {1{$random}};
  _T_1519 = _GEN_828[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_829 = {1{$random}};
  _T_1522 = _GEN_829[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_830 = {1{$random}};
  _T_1525 = _GEN_830[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_831 = {1{$random}};
  _T_1528 = _GEN_831[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_832 = {1{$random}};
  _T_1531 = _GEN_832[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_833 = {1{$random}};
  _T_1534 = _GEN_833[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_834 = {1{$random}};
  _T_1537 = _GEN_834[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_835 = {1{$random}};
  _T_1540 = _GEN_835[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_836 = {1{$random}};
  _T_1565 = _GEN_836[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_837 = {1{$random}};
  _T_1568 = _GEN_837[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_838 = {1{$random}};
  _T_1571 = _GEN_838[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_839 = {1{$random}};
  _T_1574 = _GEN_839[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_840 = {1{$random}};
  _T_1577 = _GEN_840[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_841 = {1{$random}};
  _T_1580 = _GEN_841[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_842 = {1{$random}};
  _T_1583 = _GEN_842[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_843 = {1{$random}};
  _T_1586 = _GEN_843[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_844 = {1{$random}};
  _T_1589 = _GEN_844[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_845 = {1{$random}};
  _T_1592 = _GEN_845[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_846 = {1{$random}};
  _T_1595 = _GEN_846[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_847 = {1{$random}};
  _T_1598 = _GEN_847[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_848 = {1{$random}};
  _T_1601 = _GEN_848[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_849 = {1{$random}};
  _T_1604 = _GEN_849[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_850 = {1{$random}};
  _T_1607 = _GEN_850[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_851 = {1{$random}};
  _T_1610 = _GEN_851[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_852 = {1{$random}};
  _T_1635 = _GEN_852[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_853 = {1{$random}};
  _T_1638 = _GEN_853[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_854 = {1{$random}};
  _T_1641 = _GEN_854[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_855 = {1{$random}};
  _T_1644 = _GEN_855[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_856 = {1{$random}};
  _T_1647 = _GEN_856[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_857 = {1{$random}};
  _T_1650 = _GEN_857[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_858 = {1{$random}};
  _T_1653 = _GEN_858[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_859 = {1{$random}};
  _T_1656 = _GEN_859[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_860 = {1{$random}};
  _T_1659 = _GEN_860[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_861 = {1{$random}};
  _T_1662 = _GEN_861[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_862 = {1{$random}};
  _T_1665 = _GEN_862[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_863 = {1{$random}};
  _T_1668 = _GEN_863[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_864 = {1{$random}};
  _T_1671 = _GEN_864[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_865 = {1{$random}};
  _T_1674 = _GEN_865[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_866 = {1{$random}};
  _T_1677 = _GEN_866[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_867 = {1{$random}};
  _T_1680 = _GEN_867[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_868 = {1{$random}};
  _T_1705 = _GEN_868[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_869 = {1{$random}};
  _T_1708 = _GEN_869[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_870 = {1{$random}};
  _T_1711 = _GEN_870[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_871 = {1{$random}};
  _T_1714 = _GEN_871[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_872 = {1{$random}};
  _T_1717 = _GEN_872[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_873 = {1{$random}};
  _T_1720 = _GEN_873[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_874 = {1{$random}};
  _T_1723 = _GEN_874[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_875 = {1{$random}};
  _T_1726 = _GEN_875[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_876 = {1{$random}};
  _T_1729 = _GEN_876[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_877 = {1{$random}};
  _T_1732 = _GEN_877[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_878 = {1{$random}};
  _T_1735 = _GEN_878[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_879 = {1{$random}};
  _T_1738 = _GEN_879[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_880 = {1{$random}};
  _T_1741 = _GEN_880[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_881 = {1{$random}};
  _T_1744 = _GEN_881[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_882 = {1{$random}};
  _T_1747 = _GEN_882[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_883 = {1{$random}};
  _T_1750 = _GEN_883[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_884 = {1{$random}};
  _T_1775 = _GEN_884[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_885 = {1{$random}};
  _T_1778 = _GEN_885[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_886 = {1{$random}};
  _T_1781 = _GEN_886[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_887 = {1{$random}};
  _T_1784 = _GEN_887[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_888 = {1{$random}};
  _T_1787 = _GEN_888[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_889 = {1{$random}};
  _T_1790 = _GEN_889[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_890 = {1{$random}};
  _T_1793 = _GEN_890[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_891 = {1{$random}};
  _T_1796 = _GEN_891[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_892 = {1{$random}};
  _T_1799 = _GEN_892[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_893 = {1{$random}};
  _T_1802 = _GEN_893[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_894 = {1{$random}};
  _T_1805 = _GEN_894[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_895 = {1{$random}};
  _T_1808 = _GEN_895[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_896 = {1{$random}};
  _T_1811 = _GEN_896[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_897 = {1{$random}};
  _T_1814 = _GEN_897[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_898 = {1{$random}};
  _T_1817 = _GEN_898[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_899 = {1{$random}};
  _T_1820 = _GEN_899[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_900 = {1{$random}};
  _T_1881 = _GEN_900[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_901 = {1{$random}};
  _T_1884 = _GEN_901[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_902 = {1{$random}};
  _T_1887 = _GEN_902[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_903 = {1{$random}};
  _T_1890 = _GEN_903[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_904 = {1{$random}};
  _T_1893 = _GEN_904[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_905 = {1{$random}};
  _T_1896 = _GEN_905[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_906 = {1{$random}};
  _T_1899 = _GEN_906[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_907 = {1{$random}};
  _T_1902 = _GEN_907[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_908 = {1{$random}};
  _T_1905 = _GEN_908[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_909 = {1{$random}};
  _T_1908 = _GEN_909[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_910 = {1{$random}};
  _T_1911 = _GEN_910[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_911 = {1{$random}};
  _T_1914 = _GEN_911[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_912 = {1{$random}};
  _T_1917 = _GEN_912[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_913 = {1{$random}};
  _T_1920 = _GEN_913[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_914 = {1{$random}};
  _T_1923 = _GEN_914[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_915 = {1{$random}};
  _T_1926 = _GEN_915[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_916 = {1{$random}};
  _T_1951 = _GEN_916[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_917 = {1{$random}};
  _T_1954 = _GEN_917[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_918 = {1{$random}};
  _T_1957 = _GEN_918[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_919 = {1{$random}};
  _T_1960 = _GEN_919[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_920 = {1{$random}};
  _T_1963 = _GEN_920[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_921 = {1{$random}};
  _T_1966 = _GEN_921[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_922 = {1{$random}};
  _T_1969 = _GEN_922[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_923 = {1{$random}};
  _T_1972 = _GEN_923[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_924 = {1{$random}};
  _T_1975 = _GEN_924[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_925 = {1{$random}};
  _T_1978 = _GEN_925[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_926 = {1{$random}};
  _T_1981 = _GEN_926[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_927 = {1{$random}};
  _T_1984 = _GEN_927[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_928 = {1{$random}};
  _T_1987 = _GEN_928[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_929 = {1{$random}};
  _T_1990 = _GEN_929[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_930 = {1{$random}};
  _T_1993 = _GEN_930[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_931 = {1{$random}};
  _T_1996 = _GEN_931[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_932 = {1{$random}};
  _T_2021 = _GEN_932[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_933 = {1{$random}};
  _T_2024 = _GEN_933[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_934 = {1{$random}};
  _T_2027 = _GEN_934[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_935 = {1{$random}};
  _T_2030 = _GEN_935[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_936 = {1{$random}};
  _T_2033 = _GEN_936[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_937 = {1{$random}};
  _T_2036 = _GEN_937[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_938 = {1{$random}};
  _T_2039 = _GEN_938[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_939 = {1{$random}};
  _T_2042 = _GEN_939[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_940 = {1{$random}};
  _T_2045 = _GEN_940[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_941 = {1{$random}};
  _T_2048 = _GEN_941[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_942 = {1{$random}};
  _T_2051 = _GEN_942[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_943 = {1{$random}};
  _T_2054 = _GEN_943[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_944 = {1{$random}};
  _T_2057 = _GEN_944[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_945 = {1{$random}};
  _T_2060 = _GEN_945[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_946 = {1{$random}};
  _T_2063 = _GEN_946[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_947 = {1{$random}};
  _T_2066 = _GEN_947[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_948 = {1{$random}};
  _T_2091 = _GEN_948[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_949 = {1{$random}};
  _T_2094 = _GEN_949[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_950 = {1{$random}};
  _T_2097 = _GEN_950[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_951 = {1{$random}};
  _T_2100 = _GEN_951[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_952 = {1{$random}};
  _T_2103 = _GEN_952[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_953 = {1{$random}};
  _T_2106 = _GEN_953[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_954 = {1{$random}};
  _T_2109 = _GEN_954[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_955 = {1{$random}};
  _T_2112 = _GEN_955[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_956 = {1{$random}};
  _T_2115 = _GEN_956[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_957 = {1{$random}};
  _T_2118 = _GEN_957[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_958 = {1{$random}};
  _T_2121 = _GEN_958[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_959 = {1{$random}};
  _T_2124 = _GEN_959[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_960 = {1{$random}};
  _T_2127 = _GEN_960[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_961 = {1{$random}};
  _T_2130 = _GEN_961[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_962 = {1{$random}};
  _T_2133 = _GEN_962[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_963 = {1{$random}};
  _T_2136 = _GEN_963[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_964 = {1{$random}};
  _T_2161 = _GEN_964[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_965 = {1{$random}};
  _T_2164 = _GEN_965[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_966 = {1{$random}};
  _T_2167 = _GEN_966[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_967 = {1{$random}};
  _T_2170 = _GEN_967[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_968 = {1{$random}};
  _T_2173 = _GEN_968[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_969 = {1{$random}};
  _T_2176 = _GEN_969[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_970 = {1{$random}};
  _T_2179 = _GEN_970[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_971 = {1{$random}};
  _T_2182 = _GEN_971[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_972 = {1{$random}};
  _T_2185 = _GEN_972[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_973 = {1{$random}};
  _T_2188 = _GEN_973[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_974 = {1{$random}};
  _T_2191 = _GEN_974[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_975 = {1{$random}};
  _T_2194 = _GEN_975[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_976 = {1{$random}};
  _T_2197 = _GEN_976[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_977 = {1{$random}};
  _T_2200 = _GEN_977[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_978 = {1{$random}};
  _T_2203 = _GEN_978[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_979 = {1{$random}};
  _T_2206 = _GEN_979[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_980 = {1{$random}};
  _T_2231 = _GEN_980[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_981 = {1{$random}};
  _T_2234 = _GEN_981[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_982 = {1{$random}};
  _T_2237 = _GEN_982[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_983 = {1{$random}};
  _T_2240 = _GEN_983[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_984 = {1{$random}};
  _T_2243 = _GEN_984[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_985 = {1{$random}};
  _T_2246 = _GEN_985[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_986 = {1{$random}};
  _T_2249 = _GEN_986[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_987 = {1{$random}};
  _T_2252 = _GEN_987[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_988 = {1{$random}};
  _T_2255 = _GEN_988[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_989 = {1{$random}};
  _T_2258 = _GEN_989[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_990 = {1{$random}};
  _T_2261 = _GEN_990[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_991 = {1{$random}};
  _T_2264 = _GEN_991[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_992 = {1{$random}};
  _T_2267 = _GEN_992[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_993 = {1{$random}};
  _T_2270 = _GEN_993[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_994 = {1{$random}};
  _T_2273 = _GEN_994[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_995 = {1{$random}};
  _T_2276 = _GEN_995[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_996 = {1{$random}};
  _T_2301 = _GEN_996[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_997 = {1{$random}};
  _T_2304 = _GEN_997[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_998 = {1{$random}};
  _T_2307 = _GEN_998[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_999 = {1{$random}};
  _T_2310 = _GEN_999[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1000 = {1{$random}};
  _T_2313 = _GEN_1000[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1001 = {1{$random}};
  _T_2316 = _GEN_1001[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1002 = {1{$random}};
  _T_2319 = _GEN_1002[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1003 = {1{$random}};
  _T_2322 = _GEN_1003[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1004 = {1{$random}};
  _T_2325 = _GEN_1004[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1005 = {1{$random}};
  _T_2328 = _GEN_1005[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1006 = {1{$random}};
  _T_2331 = _GEN_1006[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1007 = {1{$random}};
  _T_2334 = _GEN_1007[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1008 = {1{$random}};
  _T_2337 = _GEN_1008[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1009 = {1{$random}};
  _T_2340 = _GEN_1009[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1010 = {1{$random}};
  _T_2343 = _GEN_1010[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1011 = {1{$random}};
  _T_2346 = _GEN_1011[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1012 = {1{$random}};
  _T_2371 = _GEN_1012[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1013 = {1{$random}};
  _T_2374 = _GEN_1013[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1014 = {1{$random}};
  _T_2377 = _GEN_1014[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1015 = {1{$random}};
  _T_2380 = _GEN_1015[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1016 = {1{$random}};
  _T_2383 = _GEN_1016[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1017 = {1{$random}};
  _T_2386 = _GEN_1017[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1018 = {1{$random}};
  _T_2389 = _GEN_1018[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1019 = {1{$random}};
  _T_2392 = _GEN_1019[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1020 = {1{$random}};
  _T_2395 = _GEN_1020[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1021 = {1{$random}};
  _T_2398 = _GEN_1021[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1022 = {1{$random}};
  _T_2401 = _GEN_1022[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1023 = {1{$random}};
  _T_2404 = _GEN_1023[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1024 = {1{$random}};
  _T_2407 = _GEN_1024[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1025 = {1{$random}};
  _T_2410 = _GEN_1025[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1026 = {1{$random}};
  _T_2413 = _GEN_1026[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1027 = {1{$random}};
  _T_2416 = _GEN_1027[5:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (reset) begin
      _T_93 <= -6'sh4;
    end
    if (reset) begin
      _T_96 <= -6'sh2;
    end
    if (reset) begin
      _T_99 <= -6'sh2;
    end
    if (reset) begin
      _T_102 <= 6'sh0;
    end
    if (reset) begin
      _T_105 <= -6'sh2;
    end
    if (reset) begin
      _T_108 <= 6'sh0;
    end
    if (reset) begin
      _T_111 <= 6'sh0;
    end
    if (reset) begin
      _T_114 <= 6'sh2;
    end
    if (reset) begin
      _T_117 <= -6'sh2;
    end
    if (reset) begin
      _T_120 <= 6'sh0;
    end
    if (reset) begin
      _T_123 <= 6'sh0;
    end
    if (reset) begin
      _T_126 <= 6'sh2;
    end
    if (reset) begin
      _T_129 <= 6'sh0;
    end
    if (reset) begin
      _T_132 <= 6'sh2;
    end
    if (reset) begin
      _T_135 <= 6'sh2;
    end
    if (reset) begin
      _T_138 <= 6'sh4;
    end
    if (reset) begin
      _T_163 <= -6'sh4;
    end
    if (reset) begin
      _T_166 <= -6'sh2;
    end
    if (reset) begin
      _T_169 <= -6'sh2;
    end
    if (reset) begin
      _T_172 <= 6'sh0;
    end
    if (reset) begin
      _T_175 <= -6'sh2;
    end
    if (reset) begin
      _T_178 <= 6'sh0;
    end
    if (reset) begin
      _T_181 <= 6'sh0;
    end
    if (reset) begin
      _T_184 <= 6'sh2;
    end
    if (reset) begin
      _T_187 <= -6'sh2;
    end
    if (reset) begin
      _T_190 <= 6'sh0;
    end
    if (reset) begin
      _T_193 <= 6'sh0;
    end
    if (reset) begin
      _T_196 <= 6'sh2;
    end
    if (reset) begin
      _T_199 <= 6'sh0;
    end
    if (reset) begin
      _T_202 <= 6'sh2;
    end
    if (reset) begin
      _T_205 <= 6'sh2;
    end
    if (reset) begin
      _T_208 <= 6'sh4;
    end
    if (reset) begin
      _T_233 <= -6'sh4;
    end
    if (reset) begin
      _T_236 <= -6'sh2;
    end
    if (reset) begin
      _T_239 <= -6'sh2;
    end
    if (reset) begin
      _T_242 <= 6'sh0;
    end
    if (reset) begin
      _T_245 <= -6'sh2;
    end
    if (reset) begin
      _T_248 <= 6'sh0;
    end
    if (reset) begin
      _T_251 <= 6'sh0;
    end
    if (reset) begin
      _T_254 <= 6'sh2;
    end
    if (reset) begin
      _T_257 <= -6'sh2;
    end
    if (reset) begin
      _T_260 <= 6'sh0;
    end
    if (reset) begin
      _T_263 <= 6'sh0;
    end
    if (reset) begin
      _T_266 <= 6'sh2;
    end
    if (reset) begin
      _T_269 <= 6'sh0;
    end
    if (reset) begin
      _T_272 <= 6'sh2;
    end
    if (reset) begin
      _T_275 <= 6'sh2;
    end
    if (reset) begin
      _T_278 <= 6'sh4;
    end
    if (reset) begin
      _T_303 <= -6'sh4;
    end
    if (reset) begin
      _T_306 <= -6'sh2;
    end
    if (reset) begin
      _T_309 <= -6'sh2;
    end
    if (reset) begin
      _T_312 <= 6'sh0;
    end
    if (reset) begin
      _T_315 <= -6'sh2;
    end
    if (reset) begin
      _T_318 <= 6'sh0;
    end
    if (reset) begin
      _T_321 <= 6'sh0;
    end
    if (reset) begin
      _T_324 <= 6'sh2;
    end
    if (reset) begin
      _T_327 <= -6'sh2;
    end
    if (reset) begin
      _T_330 <= 6'sh0;
    end
    if (reset) begin
      _T_333 <= 6'sh0;
    end
    if (reset) begin
      _T_336 <= 6'sh2;
    end
    if (reset) begin
      _T_339 <= 6'sh0;
    end
    if (reset) begin
      _T_342 <= 6'sh2;
    end
    if (reset) begin
      _T_345 <= 6'sh2;
    end
    if (reset) begin
      _T_348 <= 6'sh4;
    end
    if (reset) begin
      _T_373 <= -6'sh4;
    end
    if (reset) begin
      _T_376 <= -6'sh2;
    end
    if (reset) begin
      _T_379 <= -6'sh2;
    end
    if (reset) begin
      _T_382 <= 6'sh0;
    end
    if (reset) begin
      _T_385 <= -6'sh2;
    end
    if (reset) begin
      _T_388 <= 6'sh0;
    end
    if (reset) begin
      _T_391 <= 6'sh0;
    end
    if (reset) begin
      _T_394 <= 6'sh2;
    end
    if (reset) begin
      _T_397 <= -6'sh2;
    end
    if (reset) begin
      _T_400 <= 6'sh0;
    end
    if (reset) begin
      _T_403 <= 6'sh0;
    end
    if (reset) begin
      _T_406 <= 6'sh2;
    end
    if (reset) begin
      _T_409 <= 6'sh0;
    end
    if (reset) begin
      _T_412 <= 6'sh2;
    end
    if (reset) begin
      _T_415 <= 6'sh2;
    end
    if (reset) begin
      _T_418 <= 6'sh4;
    end
    if (reset) begin
      _T_443 <= -6'sh4;
    end
    if (reset) begin
      _T_446 <= -6'sh2;
    end
    if (reset) begin
      _T_449 <= -6'sh2;
    end
    if (reset) begin
      _T_452 <= 6'sh0;
    end
    if (reset) begin
      _T_455 <= -6'sh2;
    end
    if (reset) begin
      _T_458 <= 6'sh0;
    end
    if (reset) begin
      _T_461 <= 6'sh0;
    end
    if (reset) begin
      _T_464 <= 6'sh2;
    end
    if (reset) begin
      _T_467 <= -6'sh2;
    end
    if (reset) begin
      _T_470 <= 6'sh0;
    end
    if (reset) begin
      _T_473 <= 6'sh0;
    end
    if (reset) begin
      _T_476 <= 6'sh2;
    end
    if (reset) begin
      _T_479 <= 6'sh0;
    end
    if (reset) begin
      _T_482 <= 6'sh2;
    end
    if (reset) begin
      _T_485 <= 6'sh2;
    end
    if (reset) begin
      _T_488 <= 6'sh4;
    end
    if (reset) begin
      _T_513 <= -6'sh4;
    end
    if (reset) begin
      _T_516 <= -6'sh2;
    end
    if (reset) begin
      _T_519 <= -6'sh2;
    end
    if (reset) begin
      _T_522 <= 6'sh0;
    end
    if (reset) begin
      _T_525 <= -6'sh2;
    end
    if (reset) begin
      _T_528 <= 6'sh0;
    end
    if (reset) begin
      _T_531 <= 6'sh0;
    end
    if (reset) begin
      _T_534 <= 6'sh2;
    end
    if (reset) begin
      _T_537 <= -6'sh2;
    end
    if (reset) begin
      _T_540 <= 6'sh0;
    end
    if (reset) begin
      _T_543 <= 6'sh0;
    end
    if (reset) begin
      _T_546 <= 6'sh2;
    end
    if (reset) begin
      _T_549 <= 6'sh0;
    end
    if (reset) begin
      _T_552 <= 6'sh2;
    end
    if (reset) begin
      _T_555 <= 6'sh2;
    end
    if (reset) begin
      _T_558 <= 6'sh4;
    end
    if (reset) begin
      _T_583 <= -6'sh4;
    end
    if (reset) begin
      _T_586 <= -6'sh2;
    end
    if (reset) begin
      _T_589 <= -6'sh2;
    end
    if (reset) begin
      _T_592 <= 6'sh0;
    end
    if (reset) begin
      _T_595 <= -6'sh2;
    end
    if (reset) begin
      _T_598 <= 6'sh0;
    end
    if (reset) begin
      _T_601 <= 6'sh0;
    end
    if (reset) begin
      _T_604 <= 6'sh2;
    end
    if (reset) begin
      _T_607 <= -6'sh2;
    end
    if (reset) begin
      _T_610 <= 6'sh0;
    end
    if (reset) begin
      _T_613 <= 6'sh0;
    end
    if (reset) begin
      _T_616 <= 6'sh2;
    end
    if (reset) begin
      _T_619 <= 6'sh0;
    end
    if (reset) begin
      _T_622 <= 6'sh2;
    end
    if (reset) begin
      _T_625 <= 6'sh2;
    end
    if (reset) begin
      _T_628 <= 6'sh4;
    end
    if (reset) begin
      _T_689 <= -6'sh4;
    end
    if (reset) begin
      _T_692 <= -6'sh2;
    end
    if (reset) begin
      _T_695 <= -6'sh2;
    end
    if (reset) begin
      _T_698 <= 6'sh0;
    end
    if (reset) begin
      _T_701 <= -6'sh2;
    end
    if (reset) begin
      _T_704 <= 6'sh0;
    end
    if (reset) begin
      _T_707 <= 6'sh0;
    end
    if (reset) begin
      _T_710 <= 6'sh2;
    end
    if (reset) begin
      _T_713 <= -6'sh2;
    end
    if (reset) begin
      _T_716 <= 6'sh0;
    end
    if (reset) begin
      _T_719 <= 6'sh0;
    end
    if (reset) begin
      _T_722 <= 6'sh2;
    end
    if (reset) begin
      _T_725 <= 6'sh0;
    end
    if (reset) begin
      _T_728 <= 6'sh2;
    end
    if (reset) begin
      _T_731 <= 6'sh2;
    end
    if (reset) begin
      _T_734 <= 6'sh4;
    end
    if (reset) begin
      _T_759 <= -6'sh4;
    end
    if (reset) begin
      _T_762 <= -6'sh2;
    end
    if (reset) begin
      _T_765 <= -6'sh2;
    end
    if (reset) begin
      _T_768 <= 6'sh0;
    end
    if (reset) begin
      _T_771 <= -6'sh2;
    end
    if (reset) begin
      _T_774 <= 6'sh0;
    end
    if (reset) begin
      _T_777 <= 6'sh0;
    end
    if (reset) begin
      _T_780 <= 6'sh2;
    end
    if (reset) begin
      _T_783 <= -6'sh2;
    end
    if (reset) begin
      _T_786 <= 6'sh0;
    end
    if (reset) begin
      _T_789 <= 6'sh0;
    end
    if (reset) begin
      _T_792 <= 6'sh2;
    end
    if (reset) begin
      _T_795 <= 6'sh0;
    end
    if (reset) begin
      _T_798 <= 6'sh2;
    end
    if (reset) begin
      _T_801 <= 6'sh2;
    end
    if (reset) begin
      _T_804 <= 6'sh4;
    end
    if (reset) begin
      _T_829 <= -6'sh4;
    end
    if (reset) begin
      _T_832 <= -6'sh2;
    end
    if (reset) begin
      _T_835 <= -6'sh2;
    end
    if (reset) begin
      _T_838 <= 6'sh0;
    end
    if (reset) begin
      _T_841 <= -6'sh2;
    end
    if (reset) begin
      _T_844 <= 6'sh0;
    end
    if (reset) begin
      _T_847 <= 6'sh0;
    end
    if (reset) begin
      _T_850 <= 6'sh2;
    end
    if (reset) begin
      _T_853 <= -6'sh2;
    end
    if (reset) begin
      _T_856 <= 6'sh0;
    end
    if (reset) begin
      _T_859 <= 6'sh0;
    end
    if (reset) begin
      _T_862 <= 6'sh2;
    end
    if (reset) begin
      _T_865 <= 6'sh0;
    end
    if (reset) begin
      _T_868 <= 6'sh2;
    end
    if (reset) begin
      _T_871 <= 6'sh2;
    end
    if (reset) begin
      _T_874 <= 6'sh4;
    end
    if (reset) begin
      _T_899 <= -6'sh4;
    end
    if (reset) begin
      _T_902 <= -6'sh2;
    end
    if (reset) begin
      _T_905 <= -6'sh2;
    end
    if (reset) begin
      _T_908 <= 6'sh0;
    end
    if (reset) begin
      _T_911 <= -6'sh2;
    end
    if (reset) begin
      _T_914 <= 6'sh0;
    end
    if (reset) begin
      _T_917 <= 6'sh0;
    end
    if (reset) begin
      _T_920 <= 6'sh2;
    end
    if (reset) begin
      _T_923 <= -6'sh2;
    end
    if (reset) begin
      _T_926 <= 6'sh0;
    end
    if (reset) begin
      _T_929 <= 6'sh0;
    end
    if (reset) begin
      _T_932 <= 6'sh2;
    end
    if (reset) begin
      _T_935 <= 6'sh0;
    end
    if (reset) begin
      _T_938 <= 6'sh2;
    end
    if (reset) begin
      _T_941 <= 6'sh2;
    end
    if (reset) begin
      _T_944 <= 6'sh4;
    end
    if (reset) begin
      _T_969 <= -6'sh4;
    end
    if (reset) begin
      _T_972 <= -6'sh2;
    end
    if (reset) begin
      _T_975 <= -6'sh2;
    end
    if (reset) begin
      _T_978 <= 6'sh0;
    end
    if (reset) begin
      _T_981 <= -6'sh2;
    end
    if (reset) begin
      _T_984 <= 6'sh0;
    end
    if (reset) begin
      _T_987 <= 6'sh0;
    end
    if (reset) begin
      _T_990 <= 6'sh2;
    end
    if (reset) begin
      _T_993 <= -6'sh2;
    end
    if (reset) begin
      _T_996 <= 6'sh0;
    end
    if (reset) begin
      _T_999 <= 6'sh0;
    end
    if (reset) begin
      _T_1002 <= 6'sh2;
    end
    if (reset) begin
      _T_1005 <= 6'sh0;
    end
    if (reset) begin
      _T_1008 <= 6'sh2;
    end
    if (reset) begin
      _T_1011 <= 6'sh2;
    end
    if (reset) begin
      _T_1014 <= 6'sh4;
    end
    if (reset) begin
      _T_1039 <= -6'sh4;
    end
    if (reset) begin
      _T_1042 <= -6'sh2;
    end
    if (reset) begin
      _T_1045 <= -6'sh2;
    end
    if (reset) begin
      _T_1048 <= 6'sh0;
    end
    if (reset) begin
      _T_1051 <= -6'sh2;
    end
    if (reset) begin
      _T_1054 <= 6'sh0;
    end
    if (reset) begin
      _T_1057 <= 6'sh0;
    end
    if (reset) begin
      _T_1060 <= 6'sh2;
    end
    if (reset) begin
      _T_1063 <= -6'sh2;
    end
    if (reset) begin
      _T_1066 <= 6'sh0;
    end
    if (reset) begin
      _T_1069 <= 6'sh0;
    end
    if (reset) begin
      _T_1072 <= 6'sh2;
    end
    if (reset) begin
      _T_1075 <= 6'sh0;
    end
    if (reset) begin
      _T_1078 <= 6'sh2;
    end
    if (reset) begin
      _T_1081 <= 6'sh2;
    end
    if (reset) begin
      _T_1084 <= 6'sh4;
    end
    if (reset) begin
      _T_1109 <= -6'sh4;
    end
    if (reset) begin
      _T_1112 <= -6'sh2;
    end
    if (reset) begin
      _T_1115 <= -6'sh2;
    end
    if (reset) begin
      _T_1118 <= 6'sh0;
    end
    if (reset) begin
      _T_1121 <= -6'sh2;
    end
    if (reset) begin
      _T_1124 <= 6'sh0;
    end
    if (reset) begin
      _T_1127 <= 6'sh0;
    end
    if (reset) begin
      _T_1130 <= 6'sh2;
    end
    if (reset) begin
      _T_1133 <= -6'sh2;
    end
    if (reset) begin
      _T_1136 <= 6'sh0;
    end
    if (reset) begin
      _T_1139 <= 6'sh0;
    end
    if (reset) begin
      _T_1142 <= 6'sh2;
    end
    if (reset) begin
      _T_1145 <= 6'sh0;
    end
    if (reset) begin
      _T_1148 <= 6'sh2;
    end
    if (reset) begin
      _T_1151 <= 6'sh2;
    end
    if (reset) begin
      _T_1154 <= 6'sh4;
    end
    if (reset) begin
      _T_1179 <= -6'sh4;
    end
    if (reset) begin
      _T_1182 <= -6'sh2;
    end
    if (reset) begin
      _T_1185 <= -6'sh2;
    end
    if (reset) begin
      _T_1188 <= 6'sh0;
    end
    if (reset) begin
      _T_1191 <= -6'sh2;
    end
    if (reset) begin
      _T_1194 <= 6'sh0;
    end
    if (reset) begin
      _T_1197 <= 6'sh0;
    end
    if (reset) begin
      _T_1200 <= 6'sh2;
    end
    if (reset) begin
      _T_1203 <= -6'sh2;
    end
    if (reset) begin
      _T_1206 <= 6'sh0;
    end
    if (reset) begin
      _T_1209 <= 6'sh0;
    end
    if (reset) begin
      _T_1212 <= 6'sh2;
    end
    if (reset) begin
      _T_1215 <= 6'sh0;
    end
    if (reset) begin
      _T_1218 <= 6'sh2;
    end
    if (reset) begin
      _T_1221 <= 6'sh2;
    end
    if (reset) begin
      _T_1224 <= 6'sh4;
    end
    if (reset) begin
      _T_1285 <= -6'sh4;
    end
    if (reset) begin
      _T_1288 <= -6'sh2;
    end
    if (reset) begin
      _T_1291 <= -6'sh2;
    end
    if (reset) begin
      _T_1294 <= 6'sh0;
    end
    if (reset) begin
      _T_1297 <= -6'sh2;
    end
    if (reset) begin
      _T_1300 <= 6'sh0;
    end
    if (reset) begin
      _T_1303 <= 6'sh0;
    end
    if (reset) begin
      _T_1306 <= 6'sh2;
    end
    if (reset) begin
      _T_1309 <= -6'sh2;
    end
    if (reset) begin
      _T_1312 <= 6'sh0;
    end
    if (reset) begin
      _T_1315 <= 6'sh0;
    end
    if (reset) begin
      _T_1318 <= 6'sh2;
    end
    if (reset) begin
      _T_1321 <= 6'sh0;
    end
    if (reset) begin
      _T_1324 <= 6'sh2;
    end
    if (reset) begin
      _T_1327 <= 6'sh2;
    end
    if (reset) begin
      _T_1330 <= 6'sh4;
    end
    if (reset) begin
      _T_1355 <= -6'sh4;
    end
    if (reset) begin
      _T_1358 <= -6'sh2;
    end
    if (reset) begin
      _T_1361 <= -6'sh2;
    end
    if (reset) begin
      _T_1364 <= 6'sh0;
    end
    if (reset) begin
      _T_1367 <= -6'sh2;
    end
    if (reset) begin
      _T_1370 <= 6'sh0;
    end
    if (reset) begin
      _T_1373 <= 6'sh0;
    end
    if (reset) begin
      _T_1376 <= 6'sh2;
    end
    if (reset) begin
      _T_1379 <= -6'sh2;
    end
    if (reset) begin
      _T_1382 <= 6'sh0;
    end
    if (reset) begin
      _T_1385 <= 6'sh0;
    end
    if (reset) begin
      _T_1388 <= 6'sh2;
    end
    if (reset) begin
      _T_1391 <= 6'sh0;
    end
    if (reset) begin
      _T_1394 <= 6'sh2;
    end
    if (reset) begin
      _T_1397 <= 6'sh2;
    end
    if (reset) begin
      _T_1400 <= 6'sh4;
    end
    if (reset) begin
      _T_1425 <= -6'sh4;
    end
    if (reset) begin
      _T_1428 <= -6'sh2;
    end
    if (reset) begin
      _T_1431 <= -6'sh2;
    end
    if (reset) begin
      _T_1434 <= 6'sh0;
    end
    if (reset) begin
      _T_1437 <= -6'sh2;
    end
    if (reset) begin
      _T_1440 <= 6'sh0;
    end
    if (reset) begin
      _T_1443 <= 6'sh0;
    end
    if (reset) begin
      _T_1446 <= 6'sh2;
    end
    if (reset) begin
      _T_1449 <= -6'sh2;
    end
    if (reset) begin
      _T_1452 <= 6'sh0;
    end
    if (reset) begin
      _T_1455 <= 6'sh0;
    end
    if (reset) begin
      _T_1458 <= 6'sh2;
    end
    if (reset) begin
      _T_1461 <= 6'sh0;
    end
    if (reset) begin
      _T_1464 <= 6'sh2;
    end
    if (reset) begin
      _T_1467 <= 6'sh2;
    end
    if (reset) begin
      _T_1470 <= 6'sh4;
    end
    if (reset) begin
      _T_1495 <= -6'sh4;
    end
    if (reset) begin
      _T_1498 <= -6'sh2;
    end
    if (reset) begin
      _T_1501 <= -6'sh2;
    end
    if (reset) begin
      _T_1504 <= 6'sh0;
    end
    if (reset) begin
      _T_1507 <= -6'sh2;
    end
    if (reset) begin
      _T_1510 <= 6'sh0;
    end
    if (reset) begin
      _T_1513 <= 6'sh0;
    end
    if (reset) begin
      _T_1516 <= 6'sh2;
    end
    if (reset) begin
      _T_1519 <= -6'sh2;
    end
    if (reset) begin
      _T_1522 <= 6'sh0;
    end
    if (reset) begin
      _T_1525 <= 6'sh0;
    end
    if (reset) begin
      _T_1528 <= 6'sh2;
    end
    if (reset) begin
      _T_1531 <= 6'sh0;
    end
    if (reset) begin
      _T_1534 <= 6'sh2;
    end
    if (reset) begin
      _T_1537 <= 6'sh2;
    end
    if (reset) begin
      _T_1540 <= 6'sh4;
    end
    if (reset) begin
      _T_1565 <= -6'sh4;
    end
    if (reset) begin
      _T_1568 <= -6'sh2;
    end
    if (reset) begin
      _T_1571 <= -6'sh2;
    end
    if (reset) begin
      _T_1574 <= 6'sh0;
    end
    if (reset) begin
      _T_1577 <= -6'sh2;
    end
    if (reset) begin
      _T_1580 <= 6'sh0;
    end
    if (reset) begin
      _T_1583 <= 6'sh0;
    end
    if (reset) begin
      _T_1586 <= 6'sh2;
    end
    if (reset) begin
      _T_1589 <= -6'sh2;
    end
    if (reset) begin
      _T_1592 <= 6'sh0;
    end
    if (reset) begin
      _T_1595 <= 6'sh0;
    end
    if (reset) begin
      _T_1598 <= 6'sh2;
    end
    if (reset) begin
      _T_1601 <= 6'sh0;
    end
    if (reset) begin
      _T_1604 <= 6'sh2;
    end
    if (reset) begin
      _T_1607 <= 6'sh2;
    end
    if (reset) begin
      _T_1610 <= 6'sh4;
    end
    if (reset) begin
      _T_1635 <= -6'sh4;
    end
    if (reset) begin
      _T_1638 <= -6'sh2;
    end
    if (reset) begin
      _T_1641 <= -6'sh2;
    end
    if (reset) begin
      _T_1644 <= 6'sh0;
    end
    if (reset) begin
      _T_1647 <= -6'sh2;
    end
    if (reset) begin
      _T_1650 <= 6'sh0;
    end
    if (reset) begin
      _T_1653 <= 6'sh0;
    end
    if (reset) begin
      _T_1656 <= 6'sh2;
    end
    if (reset) begin
      _T_1659 <= -6'sh2;
    end
    if (reset) begin
      _T_1662 <= 6'sh0;
    end
    if (reset) begin
      _T_1665 <= 6'sh0;
    end
    if (reset) begin
      _T_1668 <= 6'sh2;
    end
    if (reset) begin
      _T_1671 <= 6'sh0;
    end
    if (reset) begin
      _T_1674 <= 6'sh2;
    end
    if (reset) begin
      _T_1677 <= 6'sh2;
    end
    if (reset) begin
      _T_1680 <= 6'sh4;
    end
    if (reset) begin
      _T_1705 <= -6'sh4;
    end
    if (reset) begin
      _T_1708 <= -6'sh2;
    end
    if (reset) begin
      _T_1711 <= -6'sh2;
    end
    if (reset) begin
      _T_1714 <= 6'sh0;
    end
    if (reset) begin
      _T_1717 <= -6'sh2;
    end
    if (reset) begin
      _T_1720 <= 6'sh0;
    end
    if (reset) begin
      _T_1723 <= 6'sh0;
    end
    if (reset) begin
      _T_1726 <= 6'sh2;
    end
    if (reset) begin
      _T_1729 <= -6'sh2;
    end
    if (reset) begin
      _T_1732 <= 6'sh0;
    end
    if (reset) begin
      _T_1735 <= 6'sh0;
    end
    if (reset) begin
      _T_1738 <= 6'sh2;
    end
    if (reset) begin
      _T_1741 <= 6'sh0;
    end
    if (reset) begin
      _T_1744 <= 6'sh2;
    end
    if (reset) begin
      _T_1747 <= 6'sh2;
    end
    if (reset) begin
      _T_1750 <= 6'sh4;
    end
    if (reset) begin
      _T_1775 <= -6'sh4;
    end
    if (reset) begin
      _T_1778 <= -6'sh2;
    end
    if (reset) begin
      _T_1781 <= -6'sh2;
    end
    if (reset) begin
      _T_1784 <= 6'sh0;
    end
    if (reset) begin
      _T_1787 <= -6'sh2;
    end
    if (reset) begin
      _T_1790 <= 6'sh0;
    end
    if (reset) begin
      _T_1793 <= 6'sh0;
    end
    if (reset) begin
      _T_1796 <= 6'sh2;
    end
    if (reset) begin
      _T_1799 <= -6'sh2;
    end
    if (reset) begin
      _T_1802 <= 6'sh0;
    end
    if (reset) begin
      _T_1805 <= 6'sh0;
    end
    if (reset) begin
      _T_1808 <= 6'sh2;
    end
    if (reset) begin
      _T_1811 <= 6'sh0;
    end
    if (reset) begin
      _T_1814 <= 6'sh2;
    end
    if (reset) begin
      _T_1817 <= 6'sh2;
    end
    if (reset) begin
      _T_1820 <= 6'sh4;
    end
    if (reset) begin
      _T_1881 <= -6'sh4;
    end
    if (reset) begin
      _T_1884 <= -6'sh2;
    end
    if (reset) begin
      _T_1887 <= -6'sh2;
    end
    if (reset) begin
      _T_1890 <= 6'sh0;
    end
    if (reset) begin
      _T_1893 <= -6'sh2;
    end
    if (reset) begin
      _T_1896 <= 6'sh0;
    end
    if (reset) begin
      _T_1899 <= 6'sh0;
    end
    if (reset) begin
      _T_1902 <= 6'sh2;
    end
    if (reset) begin
      _T_1905 <= -6'sh2;
    end
    if (reset) begin
      _T_1908 <= 6'sh0;
    end
    if (reset) begin
      _T_1911 <= 6'sh0;
    end
    if (reset) begin
      _T_1914 <= 6'sh2;
    end
    if (reset) begin
      _T_1917 <= 6'sh0;
    end
    if (reset) begin
      _T_1920 <= 6'sh2;
    end
    if (reset) begin
      _T_1923 <= 6'sh2;
    end
    if (reset) begin
      _T_1926 <= 6'sh4;
    end
    if (reset) begin
      _T_1951 <= -6'sh4;
    end
    if (reset) begin
      _T_1954 <= -6'sh2;
    end
    if (reset) begin
      _T_1957 <= -6'sh2;
    end
    if (reset) begin
      _T_1960 <= 6'sh0;
    end
    if (reset) begin
      _T_1963 <= -6'sh2;
    end
    if (reset) begin
      _T_1966 <= 6'sh0;
    end
    if (reset) begin
      _T_1969 <= 6'sh0;
    end
    if (reset) begin
      _T_1972 <= 6'sh2;
    end
    if (reset) begin
      _T_1975 <= -6'sh2;
    end
    if (reset) begin
      _T_1978 <= 6'sh0;
    end
    if (reset) begin
      _T_1981 <= 6'sh0;
    end
    if (reset) begin
      _T_1984 <= 6'sh2;
    end
    if (reset) begin
      _T_1987 <= 6'sh0;
    end
    if (reset) begin
      _T_1990 <= 6'sh2;
    end
    if (reset) begin
      _T_1993 <= 6'sh2;
    end
    if (reset) begin
      _T_1996 <= 6'sh4;
    end
    if (reset) begin
      _T_2021 <= -6'sh4;
    end
    if (reset) begin
      _T_2024 <= -6'sh2;
    end
    if (reset) begin
      _T_2027 <= -6'sh2;
    end
    if (reset) begin
      _T_2030 <= 6'sh0;
    end
    if (reset) begin
      _T_2033 <= -6'sh2;
    end
    if (reset) begin
      _T_2036 <= 6'sh0;
    end
    if (reset) begin
      _T_2039 <= 6'sh0;
    end
    if (reset) begin
      _T_2042 <= 6'sh2;
    end
    if (reset) begin
      _T_2045 <= -6'sh2;
    end
    if (reset) begin
      _T_2048 <= 6'sh0;
    end
    if (reset) begin
      _T_2051 <= 6'sh0;
    end
    if (reset) begin
      _T_2054 <= 6'sh2;
    end
    if (reset) begin
      _T_2057 <= 6'sh0;
    end
    if (reset) begin
      _T_2060 <= 6'sh2;
    end
    if (reset) begin
      _T_2063 <= 6'sh2;
    end
    if (reset) begin
      _T_2066 <= 6'sh4;
    end
    if (reset) begin
      _T_2091 <= -6'sh4;
    end
    if (reset) begin
      _T_2094 <= -6'sh2;
    end
    if (reset) begin
      _T_2097 <= -6'sh2;
    end
    if (reset) begin
      _T_2100 <= 6'sh0;
    end
    if (reset) begin
      _T_2103 <= -6'sh2;
    end
    if (reset) begin
      _T_2106 <= 6'sh0;
    end
    if (reset) begin
      _T_2109 <= 6'sh0;
    end
    if (reset) begin
      _T_2112 <= 6'sh2;
    end
    if (reset) begin
      _T_2115 <= -6'sh2;
    end
    if (reset) begin
      _T_2118 <= 6'sh0;
    end
    if (reset) begin
      _T_2121 <= 6'sh0;
    end
    if (reset) begin
      _T_2124 <= 6'sh2;
    end
    if (reset) begin
      _T_2127 <= 6'sh0;
    end
    if (reset) begin
      _T_2130 <= 6'sh2;
    end
    if (reset) begin
      _T_2133 <= 6'sh2;
    end
    if (reset) begin
      _T_2136 <= 6'sh4;
    end
    if (reset) begin
      _T_2161 <= -6'sh4;
    end
    if (reset) begin
      _T_2164 <= -6'sh2;
    end
    if (reset) begin
      _T_2167 <= -6'sh2;
    end
    if (reset) begin
      _T_2170 <= 6'sh0;
    end
    if (reset) begin
      _T_2173 <= -6'sh2;
    end
    if (reset) begin
      _T_2176 <= 6'sh0;
    end
    if (reset) begin
      _T_2179 <= 6'sh0;
    end
    if (reset) begin
      _T_2182 <= 6'sh2;
    end
    if (reset) begin
      _T_2185 <= -6'sh2;
    end
    if (reset) begin
      _T_2188 <= 6'sh0;
    end
    if (reset) begin
      _T_2191 <= 6'sh0;
    end
    if (reset) begin
      _T_2194 <= 6'sh2;
    end
    if (reset) begin
      _T_2197 <= 6'sh0;
    end
    if (reset) begin
      _T_2200 <= 6'sh2;
    end
    if (reset) begin
      _T_2203 <= 6'sh2;
    end
    if (reset) begin
      _T_2206 <= 6'sh4;
    end
    if (reset) begin
      _T_2231 <= -6'sh4;
    end
    if (reset) begin
      _T_2234 <= -6'sh2;
    end
    if (reset) begin
      _T_2237 <= -6'sh2;
    end
    if (reset) begin
      _T_2240 <= 6'sh0;
    end
    if (reset) begin
      _T_2243 <= -6'sh2;
    end
    if (reset) begin
      _T_2246 <= 6'sh0;
    end
    if (reset) begin
      _T_2249 <= 6'sh0;
    end
    if (reset) begin
      _T_2252 <= 6'sh2;
    end
    if (reset) begin
      _T_2255 <= -6'sh2;
    end
    if (reset) begin
      _T_2258 <= 6'sh0;
    end
    if (reset) begin
      _T_2261 <= 6'sh0;
    end
    if (reset) begin
      _T_2264 <= 6'sh2;
    end
    if (reset) begin
      _T_2267 <= 6'sh0;
    end
    if (reset) begin
      _T_2270 <= 6'sh2;
    end
    if (reset) begin
      _T_2273 <= 6'sh2;
    end
    if (reset) begin
      _T_2276 <= 6'sh4;
    end
    if (reset) begin
      _T_2301 <= -6'sh4;
    end
    if (reset) begin
      _T_2304 <= -6'sh2;
    end
    if (reset) begin
      _T_2307 <= -6'sh2;
    end
    if (reset) begin
      _T_2310 <= 6'sh0;
    end
    if (reset) begin
      _T_2313 <= -6'sh2;
    end
    if (reset) begin
      _T_2316 <= 6'sh0;
    end
    if (reset) begin
      _T_2319 <= 6'sh0;
    end
    if (reset) begin
      _T_2322 <= 6'sh2;
    end
    if (reset) begin
      _T_2325 <= -6'sh2;
    end
    if (reset) begin
      _T_2328 <= 6'sh0;
    end
    if (reset) begin
      _T_2331 <= 6'sh0;
    end
    if (reset) begin
      _T_2334 <= 6'sh2;
    end
    if (reset) begin
      _T_2337 <= 6'sh0;
    end
    if (reset) begin
      _T_2340 <= 6'sh2;
    end
    if (reset) begin
      _T_2343 <= 6'sh2;
    end
    if (reset) begin
      _T_2346 <= 6'sh4;
    end
    if (reset) begin
      _T_2371 <= -6'sh4;
    end
    if (reset) begin
      _T_2374 <= -6'sh2;
    end
    if (reset) begin
      _T_2377 <= -6'sh2;
    end
    if (reset) begin
      _T_2380 <= 6'sh0;
    end
    if (reset) begin
      _T_2383 <= -6'sh2;
    end
    if (reset) begin
      _T_2386 <= 6'sh0;
    end
    if (reset) begin
      _T_2389 <= 6'sh0;
    end
    if (reset) begin
      _T_2392 <= 6'sh2;
    end
    if (reset) begin
      _T_2395 <= -6'sh2;
    end
    if (reset) begin
      _T_2398 <= 6'sh0;
    end
    if (reset) begin
      _T_2401 <= 6'sh0;
    end
    if (reset) begin
      _T_2404 <= 6'sh2;
    end
    if (reset) begin
      _T_2407 <= 6'sh0;
    end
    if (reset) begin
      _T_2410 <= 6'sh2;
    end
    if (reset) begin
      _T_2413 <= 6'sh2;
    end
    if (reset) begin
      _T_2416 <= 6'sh4;
    end
  end
endmodule
module IglooScheduler(
  input        clock,
  input        reset,
  input        io_en,
  input  [7:0] io_inputOffset,
  input  [7:0] io_memOffset,
  output       io_finished,
  output [3:0] io_result
);
  wire  hw_clock;
  wire  hw_reset;
  wire [3:0] hw_io_input;
  wire  hw_io_inputSel;
  wire  hw_io_inputBufferPush;
  wire  hw_io_inputBufferPop;
  wire  hw_io_memSel;
  wire [7:0] hw_io_memAddr;
  wire [127:0] hw_io_memOut;
  wire  hw_io_memRen;
  wire  hw_io_memWen;
  wire [127:0] hw_io_memIn;
  wire  hw_io_accEn;
  wire [4:0] hw_io_accSel;
  wire  hw_io_accReset;
  wire  hw_io_maxClear;
  wire  hw_io_maxEn;
  wire [3:0] hw_io_maxOffset;
  wire  hw_io_meanReset;
  wire [15:0] hw_io_featureNumInverse65536;
  wire  hw_io_meanUpdate;
  wire [3:0] hw_io_result;
  reg [3:0] currentLayer;
  reg [31:0] _GEN_45;
  wire  _T_15;
  wire [3:0] _T_16;
  wire  _T_17;
  wire [6:0] currentFeatureCnt;
  wire [6:0] accWidth;
  wire [1:0] _T_25;
  wire [3:0] inputRound;
  wire [6:0] _GEN_158;
  wire [10:0] currentTotalRound;
  wire  _T_28;
  reg [7:0] state;
  reg [31:0] _GEN_46;
  reg [15:0] substate;
  reg [31:0] _GEN_47;
  wire [127:0] _T_35;
  wire [3:0] inputBuffer_0;
  wire [3:0] inputBuffer_1;
  wire [3:0] inputBuffer_2;
  wire [3:0] inputBuffer_3;
  wire [3:0] inputBuffer_4;
  wire [3:0] inputBuffer_5;
  wire [3:0] inputBuffer_6;
  wire [3:0] inputBuffer_7;
  wire [3:0] inputBuffer_8;
  wire [3:0] inputBuffer_9;
  wire [3:0] inputBuffer_10;
  wire [3:0] inputBuffer_11;
  wire [3:0] inputBuffer_12;
  wire [3:0] inputBuffer_13;
  wire [3:0] inputBuffer_14;
  wire [3:0] inputBuffer_15;
  wire [3:0] inputBuffer_16;
  wire [3:0] inputBuffer_17;
  wire [3:0] inputBuffer_18;
  wire [3:0] inputBuffer_19;
  wire [3:0] inputBuffer_20;
  wire [3:0] inputBuffer_21;
  wire [3:0] inputBuffer_22;
  wire [3:0] inputBuffer_23;
  wire [3:0] inputBuffer_24;
  wire [3:0] inputBuffer_25;
  wire [3:0] inputBuffer_26;
  wire [3:0] inputBuffer_27;
  wire [3:0] inputBuffer_28;
  wire [3:0] inputBuffer_29;
  wire [3:0] inputBuffer_30;
  wire [3:0] inputBuffer_31;
  wire [127:0] _T_142;
  wire [3:0] _T_143;
  wire [3:0] _T_144;
  wire [3:0] _T_145;
  wire [3:0] _T_146;
  wire [3:0] _T_147;
  wire [3:0] _T_148;
  wire [3:0] _T_149;
  wire [3:0] _T_150;
  wire [3:0] _T_151;
  wire [3:0] _T_152;
  wire [3:0] _T_153;
  wire [3:0] _T_154;
  wire [3:0] _T_155;
  wire [3:0] _T_156;
  wire [3:0] _T_157;
  wire [3:0] _T_158;
  wire [3:0] _T_159;
  wire [3:0] _T_160;
  wire [3:0] _T_161;
  wire [3:0] _T_162;
  wire [3:0] _T_163;
  wire [3:0] _T_164;
  wire [3:0] _T_165;
  wire [3:0] _T_166;
  wire [3:0] _T_167;
  wire [3:0] _T_168;
  wire [3:0] _T_169;
  wire [3:0] _T_170;
  wire [3:0] _T_171;
  wire [3:0] _T_172;
  wire [3:0] _T_173;
  wire [3:0] _T_174;
  reg [3:0] maxOffsetReg;
  reg [31:0] _GEN_48;
  wire  _T_177;
  wire [3:0] _GEN_4;
  wire [7:0] _GEN_5;
  wire [15:0] _GEN_6;
  wire  _T_186;
  wire [7:0] _GEN_7;
  wire [15:0] _GEN_8;
  wire  _T_190;
  wire  _T_194;
  wire [16:0] _T_196;
  wire [16:0] _T_197;
  wire [15:0] _T_198;
  wire [4:0] _T_201;
  wire [3:0] _GEN_0;
  wire [3:0] _GEN_9;
  wire [3:0] _GEN_10;
  wire [3:0] _GEN_11;
  wire [3:0] _GEN_12;
  wire [3:0] _GEN_13;
  wire [3:0] _GEN_14;
  wire [3:0] _GEN_15;
  wire [3:0] _GEN_16;
  wire [3:0] _GEN_17;
  wire [3:0] _GEN_18;
  wire [3:0] _GEN_19;
  wire [3:0] _GEN_20;
  wire [3:0] _GEN_21;
  wire [3:0] _GEN_22;
  wire [3:0] _GEN_23;
  wire [3:0] _GEN_24;
  wire [3:0] _GEN_25;
  wire [3:0] _GEN_26;
  wire [3:0] _GEN_27;
  wire [3:0] _GEN_28;
  wire [3:0] _GEN_29;
  wire [3:0] _GEN_30;
  wire [3:0] _GEN_31;
  wire [3:0] _GEN_32;
  wire [3:0] _GEN_33;
  wire [3:0] _GEN_34;
  wire [3:0] _GEN_35;
  wire [3:0] _GEN_36;
  wire [3:0] _GEN_37;
  wire [3:0] _GEN_38;
  wire [3:0] _GEN_39;
  wire [16:0] _T_203;
  wire [15:0] _T_204;
  wire [15:0] _GEN_41;
  wire  _T_206;
  wire  _T_208;
  wire  _T_209;
  wire [3:0] _GEN_1;
  wire [3:0] _GEN_73;
  wire [7:0] _GEN_74;
  wire [7:0] _GEN_75;
  wire [15:0] _GEN_76;
  wire [15:0] _GEN_80;
  wire [7:0] _GEN_81;
  wire [7:0] _GEN_82;
  wire  _T_220;
  wire [8:0] _T_226;
  wire [7:0] _T_227;
  wire  _GEN_83;
  wire [7:0] _GEN_87;
  wire [7:0] _GEN_88;
  wire [15:0] _GEN_89;
  wire  _T_231;
  wire [15:0] _GEN_159;
  wire [15:0] _GEN_2;
  wire [6:0] _T_235;
  wire [15:0] _GEN_160;
  wire [16:0] _T_236;
  wire [15:0] _T_237;
  wire [16:0] _T_239;
  wire [15:0] _T_240;
  wire [11:0] _T_242;
  wire [11:0] _T_243;
  wire [10:0] _T_244;
  wire [15:0] _GEN_161;
  wire  _T_245;
  wire [15:0] _GEN_90;
  wire  _T_253;
  wire  _T_255;
  wire  _T_256;
  wire  _GEN_91;
  wire  _GEN_92;
  wire [7:0] _GEN_93;
  wire [15:0] _GEN_94;
  wire [3:0] _GEN_96;
  wire [15:0] _GEN_3;
  wire [6:0] _T_263;
  wire [7:0] _T_265;
  wire [7:0] _T_266;
  wire [6:0] _T_267;
  wire  _T_268;
  wire [7:0] _T_272;
  wire [7:0] _T_273;
  wire [6:0] _T_274;
  wire  _T_275;
  wire  _T_277;
  wire  _T_278;
  wire  _GEN_99;
  wire [6:0] _GEN_100;
  wire [15:0] _GEN_101;
  wire [15:0] _GEN_102;
  wire  _GEN_103;
  wire  _GEN_104;
  wire [7:0] _GEN_105;
  wire [3:0] _GEN_107;
  wire  _GEN_109;
  wire  _T_281;
  wire [15:0] _GEN_165;
  wire  _T_286;
  wire  _GEN_111;
  wire [7:0] _GEN_112;
  wire  _T_292;
  wire [4:0] _T_294;
  wire [3:0] _T_295;
  wire [3:0] _GEN_114;
  wire  _GEN_115;
  wire  _GEN_117;
  wire [7:0] _GEN_119;
  wire  _GEN_122;
  wire [7:0] _GEN_123;
  wire [3:0] _GEN_125;
  wire  _GEN_126;
  wire  _GEN_128;
  wire [15:0] _GEN_167;
  wire [16:0] _T_307;
  wire [15:0] _T_308;
  wire [16:0] _T_310;
  wire [15:0] _T_311;
  wire [4:0] _T_314;
  wire [3:0] _T_315;
  wire  _GEN_131;
  wire [7:0] _GEN_132;
  wire [15:0] _GEN_133;
  wire [3:0] _GEN_134;
  wire  _GEN_135;
  wire  _GEN_137;
  wire [15:0] _GEN_138;
  wire [15:0] _GEN_139;
  wire  _GEN_140;
  wire [3:0] _GEN_141;
  wire [3:0] _GEN_145;
  wire [7:0] _GEN_146;
  wire [15:0] _GEN_147;
  wire [3:0] _GEN_155;
  wire  _GEN_157;
  reg [127:0] _GEN_40;
  reg [127:0] _GEN_49;
  reg  _GEN_42;
  reg [31:0] _GEN_50;
  reg [15:0] _GEN_43;
  reg [31:0] _GEN_51;
  reg  _GEN_44;
  reg [31:0] _GEN_52;
  XNORNetInference hw (
    .clock(hw_clock),
    .reset(hw_reset),
    .io_input(hw_io_input),
    .io_inputSel(hw_io_inputSel),
    .io_inputBufferPush(hw_io_inputBufferPush),
    .io_inputBufferPop(hw_io_inputBufferPop),
    .io_memSel(hw_io_memSel),
    .io_memAddr(hw_io_memAddr),
    .io_memOut(hw_io_memOut),
    .io_memRen(hw_io_memRen),
    .io_memWen(hw_io_memWen),
    .io_memIn(hw_io_memIn),
    .io_accEn(hw_io_accEn),
    .io_accSel(hw_io_accSel),
    .io_accReset(hw_io_accReset),
    .io_maxClear(hw_io_maxClear),
    .io_maxEn(hw_io_maxEn),
    .io_maxOffset(hw_io_maxOffset),
    .io_meanReset(hw_io_meanReset),
    .io_featureNumInverse65536(hw_io_featureNumInverse65536),
    .io_meanUpdate(hw_io_meanUpdate),
    .io_result(hw_io_result)
  );
  assign io_finished = 1'h1;
  assign io_result = hw_io_result;
  assign hw_clock = clock;
  assign hw_reset = reset;
  assign hw_io_input = _GEN_73;
  assign hw_io_inputSel = _GEN_83;
  assign hw_io_inputBufferPush = _GEN_135;
  assign hw_io_inputBufferPop = _GEN_109;
  assign hw_io_memSel = _GEN_103;
  assign hw_io_memAddr = _GEN_139[7:0];
  assign hw_io_memRen = 1'h1;
  assign hw_io_memWen = 1'h0;
  assign hw_io_memIn = _GEN_40;
  assign hw_io_accEn = _GEN_137;
  assign hw_io_accSel = _GEN_138[4:0];
  assign hw_io_accReset = 1'h1;
  assign hw_io_maxClear = _GEN_140;
  assign hw_io_maxEn = _GEN_157;
  assign hw_io_maxOffset = maxOffsetReg;
  assign hw_io_meanReset = _GEN_42;
  assign hw_io_featureNumInverse65536 = _GEN_43;
  assign hw_io_meanUpdate = _GEN_44;
  assign _T_15 = 4'h1 == currentLayer;
  assign _T_16 = _T_15 ? 4'hc : 4'h0;
  assign _T_17 = 4'h0 == currentLayer;
  assign currentFeatureCnt = _T_17 ? 7'h60 : {{3'd0}, _T_16};
  assign accWidth = currentFeatureCnt / 7'h4;
  assign _T_25 = _T_15 ? 2'h3 : 2'h0;
  assign inputRound = _T_17 ? 4'h8 : {{2'd0}, _T_25};
  assign _GEN_158 = {{3'd0}, inputRound};
  assign currentTotalRound = accWidth * _GEN_158;
  assign _T_28 = currentLayer == 4'h1;
  assign _T_35 = hw_io_memOut;
  assign inputBuffer_0 = _T_143;
  assign inputBuffer_1 = _T_144;
  assign inputBuffer_2 = _T_145;
  assign inputBuffer_3 = _T_146;
  assign inputBuffer_4 = _T_147;
  assign inputBuffer_5 = _T_148;
  assign inputBuffer_6 = _T_149;
  assign inputBuffer_7 = _T_150;
  assign inputBuffer_8 = _T_151;
  assign inputBuffer_9 = _T_152;
  assign inputBuffer_10 = _T_153;
  assign inputBuffer_11 = _T_154;
  assign inputBuffer_12 = _T_155;
  assign inputBuffer_13 = _T_156;
  assign inputBuffer_14 = _T_157;
  assign inputBuffer_15 = _T_158;
  assign inputBuffer_16 = _T_159;
  assign inputBuffer_17 = _T_160;
  assign inputBuffer_18 = _T_161;
  assign inputBuffer_19 = _T_162;
  assign inputBuffer_20 = _T_163;
  assign inputBuffer_21 = _T_164;
  assign inputBuffer_22 = _T_165;
  assign inputBuffer_23 = _T_166;
  assign inputBuffer_24 = _T_167;
  assign inputBuffer_25 = _T_168;
  assign inputBuffer_26 = _T_169;
  assign inputBuffer_27 = _T_170;
  assign inputBuffer_28 = _T_171;
  assign inputBuffer_29 = _T_172;
  assign inputBuffer_30 = _T_173;
  assign inputBuffer_31 = _T_174;
  assign _T_142 = _T_35;
  assign _T_143 = _T_142[3:0];
  assign _T_144 = _T_142[7:4];
  assign _T_145 = _T_142[11:8];
  assign _T_146 = _T_142[15:12];
  assign _T_147 = _T_142[19:16];
  assign _T_148 = _T_142[23:20];
  assign _T_149 = _T_142[27:24];
  assign _T_150 = _T_142[31:28];
  assign _T_151 = _T_142[35:32];
  assign _T_152 = _T_142[39:36];
  assign _T_153 = _T_142[43:40];
  assign _T_154 = _T_142[47:44];
  assign _T_155 = _T_142[51:48];
  assign _T_156 = _T_142[55:52];
  assign _T_157 = _T_142[59:56];
  assign _T_158 = _T_142[63:60];
  assign _T_159 = _T_142[67:64];
  assign _T_160 = _T_142[71:68];
  assign _T_161 = _T_142[75:72];
  assign _T_162 = _T_142[79:76];
  assign _T_163 = _T_142[83:80];
  assign _T_164 = _T_142[87:84];
  assign _T_165 = _T_142[91:88];
  assign _T_166 = _T_142[95:92];
  assign _T_167 = _T_142[99:96];
  assign _T_168 = _T_142[103:100];
  assign _T_169 = _T_142[107:104];
  assign _T_170 = _T_142[111:108];
  assign _T_171 = _T_142[115:112];
  assign _T_172 = _T_142[119:116];
  assign _T_173 = _T_142[123:120];
  assign _T_174 = _T_142[127:124];
  assign _T_177 = state == 8'h0;
  assign _GEN_4 = _T_177 ? 4'h0 : currentLayer;
  assign _GEN_5 = _T_177 ? 8'h1 : state;
  assign _GEN_6 = _T_177 ? 16'h0 : substate;
  assign _T_186 = state == 8'h1;
  assign _GEN_7 = _T_186 ? 8'h2 : _GEN_5;
  assign _GEN_8 = _T_186 ? 16'h0 : _GEN_6;
  assign _T_190 = state == 8'h2;
  assign _T_194 = substate < 16'h1f;
  assign _T_196 = 16'h1f - substate;
  assign _T_197 = $unsigned(_T_196);
  assign _T_198 = _T_197[15:0];
  assign _T_201 = _T_198[4:0];
  assign _GEN_0 = _GEN_39;
  assign _GEN_9 = 5'h1 == _T_201 ? inputBuffer_1 : inputBuffer_0;
  assign _GEN_10 = 5'h2 == _T_201 ? inputBuffer_2 : _GEN_9;
  assign _GEN_11 = 5'h3 == _T_201 ? inputBuffer_3 : _GEN_10;
  assign _GEN_12 = 5'h4 == _T_201 ? inputBuffer_4 : _GEN_11;
  assign _GEN_13 = 5'h5 == _T_201 ? inputBuffer_5 : _GEN_12;
  assign _GEN_14 = 5'h6 == _T_201 ? inputBuffer_6 : _GEN_13;
  assign _GEN_15 = 5'h7 == _T_201 ? inputBuffer_7 : _GEN_14;
  assign _GEN_16 = 5'h8 == _T_201 ? inputBuffer_8 : _GEN_15;
  assign _GEN_17 = 5'h9 == _T_201 ? inputBuffer_9 : _GEN_16;
  assign _GEN_18 = 5'ha == _T_201 ? inputBuffer_10 : _GEN_17;
  assign _GEN_19 = 5'hb == _T_201 ? inputBuffer_11 : _GEN_18;
  assign _GEN_20 = 5'hc == _T_201 ? inputBuffer_12 : _GEN_19;
  assign _GEN_21 = 5'hd == _T_201 ? inputBuffer_13 : _GEN_20;
  assign _GEN_22 = 5'he == _T_201 ? inputBuffer_14 : _GEN_21;
  assign _GEN_23 = 5'hf == _T_201 ? inputBuffer_15 : _GEN_22;
  assign _GEN_24 = 5'h10 == _T_201 ? inputBuffer_16 : _GEN_23;
  assign _GEN_25 = 5'h11 == _T_201 ? inputBuffer_17 : _GEN_24;
  assign _GEN_26 = 5'h12 == _T_201 ? inputBuffer_18 : _GEN_25;
  assign _GEN_27 = 5'h13 == _T_201 ? inputBuffer_19 : _GEN_26;
  assign _GEN_28 = 5'h14 == _T_201 ? inputBuffer_20 : _GEN_27;
  assign _GEN_29 = 5'h15 == _T_201 ? inputBuffer_21 : _GEN_28;
  assign _GEN_30 = 5'h16 == _T_201 ? inputBuffer_22 : _GEN_29;
  assign _GEN_31 = 5'h17 == _T_201 ? inputBuffer_23 : _GEN_30;
  assign _GEN_32 = 5'h18 == _T_201 ? inputBuffer_24 : _GEN_31;
  assign _GEN_33 = 5'h19 == _T_201 ? inputBuffer_25 : _GEN_32;
  assign _GEN_34 = 5'h1a == _T_201 ? inputBuffer_26 : _GEN_33;
  assign _GEN_35 = 5'h1b == _T_201 ? inputBuffer_27 : _GEN_34;
  assign _GEN_36 = 5'h1c == _T_201 ? inputBuffer_28 : _GEN_35;
  assign _GEN_37 = 5'h1d == _T_201 ? inputBuffer_29 : _GEN_36;
  assign _GEN_38 = 5'h1e == _T_201 ? inputBuffer_30 : _GEN_37;
  assign _GEN_39 = 5'h1f == _T_201 ? inputBuffer_31 : _GEN_38;
  assign _T_203 = substate + 16'h1;
  assign _T_204 = _T_203[15:0];
  assign _GEN_41 = _T_194 ? _T_204 : _GEN_8;
  assign _T_206 = substate == 16'h1f;
  assign _T_208 = _T_194 == 1'h0;
  assign _T_209 = _T_208 & _T_206;
  assign _GEN_1 = _GEN_39;
  assign _GEN_73 = _T_209 ? _GEN_1 : _GEN_0;
  assign _GEN_74 = _T_209 ? io_memOffset : io_inputOffset;
  assign _GEN_75 = _T_209 ? 8'h3 : _GEN_7;
  assign _GEN_76 = _T_209 ? 16'h0 : _GEN_41;
  assign _GEN_80 = _T_190 ? _GEN_76 : _GEN_8;
  assign _GEN_81 = _T_190 ? _GEN_74 : io_inputOffset;
  assign _GEN_82 = _T_190 ? _GEN_75 : _GEN_7;
  assign _T_220 = state == 8'h3;
  assign _T_226 = io_memOffset + 8'h1;
  assign _T_227 = _T_226[7:0];
  assign _GEN_83 = _T_220 ? 1'h0 : 1'h1;
  assign _GEN_87 = _T_220 ? _T_227 : _GEN_81;
  assign _GEN_88 = _T_220 ? 8'h4 : _GEN_82;
  assign _GEN_89 = _T_220 ? 16'h0 : _GEN_80;
  assign _T_231 = state == 8'h4;
  assign _GEN_159 = {{9'd0}, accWidth};
  assign _GEN_2 = _T_204 % _GEN_159;
  assign _T_235 = _GEN_2[6:0];
  assign _GEN_160 = {{8'd0}, io_memOffset};
  assign _T_236 = _GEN_160 + substate;
  assign _T_237 = _T_236[15:0];
  assign _T_239 = _T_237 + 16'h2;
  assign _T_240 = _T_239[15:0];
  assign _T_242 = currentTotalRound - 11'h1;
  assign _T_243 = $unsigned(_T_242);
  assign _T_244 = _T_243[10:0];
  assign _GEN_161 = {{5'd0}, _T_244};
  assign _T_245 = substate < _GEN_161;
  assign _GEN_90 = _T_245 ? _T_204 : _GEN_89;
  assign _T_253 = substate == _GEN_161;
  assign _T_255 = _T_245 == 1'h0;
  assign _T_256 = _T_255 & _T_253;
  assign _GEN_91 = _T_256 ? 1'h0 : 1'h1;
  assign _GEN_92 = _T_256 ? 1'h1 : _GEN_83;
  assign _GEN_93 = _T_256 ? 8'h5 : _GEN_88;
  assign _GEN_94 = _T_256 ? 16'h0 : _GEN_90;
  assign _GEN_96 = _T_256 ? 4'h0 : maxOffsetReg;
  assign _GEN_3 = substate % _GEN_159;
  assign _T_263 = _GEN_3[6:0];
  assign _T_265 = accWidth - 7'h2;
  assign _T_266 = $unsigned(_T_265);
  assign _T_267 = _T_266[6:0];
  assign _T_268 = _T_263 == _T_267;
  assign _T_272 = accWidth - 7'h1;
  assign _T_273 = $unsigned(_T_272);
  assign _T_274 = _T_273[6:0];
  assign _T_275 = _T_263 == _T_274;
  assign _T_277 = _T_268 == 1'h0;
  assign _T_278 = _T_277 & _T_275;
  assign _GEN_99 = _T_278 ? 1'h0 : _T_268;
  assign _GEN_100 = _T_231 ? _T_235 : 7'h0;
  assign _GEN_101 = _T_231 ? _T_240 : {{8'd0}, _GEN_87};
  assign _GEN_102 = _T_231 ? _GEN_94 : _GEN_89;
  assign _GEN_103 = _T_231 ? _GEN_91 : 1'h1;
  assign _GEN_104 = _T_231 ? _GEN_92 : _GEN_83;
  assign _GEN_105 = _T_231 ? _GEN_93 : _GEN_88;
  assign _GEN_107 = _T_231 ? _GEN_96 : maxOffsetReg;
  assign _GEN_109 = _T_231 ? _GEN_99 : 1'h0;
  assign _T_281 = state == 8'h5;
  assign _GEN_165 = {{9'd0}, _T_274};
  assign _T_286 = substate == _GEN_165;
  assign _GEN_111 = _T_28 ? 1'h0 : _T_28;
  assign _GEN_112 = _T_28 ? 8'h6 : _GEN_105;
  assign _T_292 = _T_28 == 1'h0;
  assign _T_294 = currentLayer + 4'h1;
  assign _T_295 = _T_294[3:0];
  assign _GEN_114 = _T_292 ? _T_295 : _GEN_4;
  assign _GEN_115 = _T_292 ? 1'h0 : _GEN_104;
  assign _GEN_117 = _T_292 ? 1'h1 : _GEN_103;
  assign _GEN_119 = _T_292 ? 8'h4 : _GEN_112;
  assign _GEN_122 = _T_286 ? _GEN_111 : _T_28;
  assign _GEN_123 = _T_286 ? _GEN_119 : _GEN_105;
  assign _GEN_125 = _T_286 ? _GEN_114 : _GEN_4;
  assign _GEN_126 = _T_286 ? _GEN_115 : _GEN_104;
  assign _GEN_128 = _T_286 ? _GEN_117 : _GEN_103;
  assign _GEN_167 = {{5'd0}, currentTotalRound};
  assign _T_307 = _T_237 + _GEN_167;
  assign _T_308 = _T_307[15:0];
  assign _T_310 = _T_308 + 16'h2;
  assign _T_311 = _T_310[15:0];
  assign _T_314 = maxOffsetReg + 4'h4;
  assign _T_315 = _T_314[3:0];
  assign _GEN_131 = _T_281 ? _GEN_122 : _T_28;
  assign _GEN_132 = _T_281 ? _GEN_123 : _GEN_105;
  assign _GEN_133 = _T_281 ? _T_204 : _GEN_102;
  assign _GEN_134 = _T_281 ? _GEN_125 : _GEN_4;
  assign _GEN_135 = _T_281 ? _GEN_126 : _GEN_104;
  assign _GEN_137 = _T_281 ? _GEN_128 : _GEN_103;
  assign _GEN_138 = _T_281 ? _T_204 : {{9'd0}, _GEN_100};
  assign _GEN_139 = _T_281 ? _T_311 : _GEN_101;
  assign _GEN_140 = _T_281 ? 1'h0 : 1'h1;
  assign _GEN_141 = _T_281 ? _T_315 : _GEN_107;
  assign _GEN_145 = io_en ? _GEN_134 : currentLayer;
  assign _GEN_146 = io_en ? _GEN_132 : state;
  assign _GEN_147 = io_en ? _GEN_133 : substate;
  assign _GEN_155 = io_en ? _GEN_141 : maxOffsetReg;
  assign _GEN_157 = io_en ? _GEN_131 : _T_28;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_45 = {1{$random}};
  currentLayer = _GEN_45[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_46 = {1{$random}};
  state = _GEN_46[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_47 = {1{$random}};
  substate = _GEN_47[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_48 = {1{$random}};
  maxOffsetReg = _GEN_48[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_49 = {4{$random}};
  _GEN_40 = _GEN_49[127:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_50 = {1{$random}};
  _GEN_42 = _GEN_50[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_51 = {1{$random}};
  _GEN_43 = _GEN_51[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_52 = {1{$random}};
  _GEN_44 = _GEN_52[0:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (io_en) begin
      if (_T_281) begin
        if (_T_286) begin
          if (_T_292) begin
            currentLayer <= _T_295;
          end else begin
            if (_T_177) begin
              currentLayer <= 4'h0;
            end
          end
        end else begin
          if (_T_177) begin
            currentLayer <= 4'h0;
          end
        end
      end else begin
        if (_T_177) begin
          currentLayer <= 4'h0;
        end
      end
    end
    if (reset) begin
      state <= 8'h0;
    end else begin
      if (io_en) begin
        if (_T_281) begin
          if (_T_286) begin
            if (_T_292) begin
              state <= 8'h4;
            end else begin
              if (_T_28) begin
                state <= 8'h6;
              end else begin
                if (_T_231) begin
                  if (_T_256) begin
                    state <= 8'h5;
                  end else begin
                    if (_T_220) begin
                      state <= 8'h4;
                    end else begin
                      if (_T_190) begin
                        if (_T_209) begin
                          state <= 8'h3;
                        end else begin
                          if (_T_186) begin
                            state <= 8'h2;
                          end else begin
                            if (_T_177) begin
                              state <= 8'h1;
                            end
                          end
                        end
                      end else begin
                        if (_T_186) begin
                          state <= 8'h2;
                        end else begin
                          if (_T_177) begin
                            state <= 8'h1;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if (_T_220) begin
                    state <= 8'h4;
                  end else begin
                    if (_T_190) begin
                      if (_T_209) begin
                        state <= 8'h3;
                      end else begin
                        if (_T_186) begin
                          state <= 8'h2;
                        end else begin
                          if (_T_177) begin
                            state <= 8'h1;
                          end
                        end
                      end
                    end else begin
                      if (_T_186) begin
                        state <= 8'h2;
                      end else begin
                        if (_T_177) begin
                          state <= 8'h1;
                        end
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_231) begin
              if (_T_256) begin
                state <= 8'h5;
              end else begin
                if (_T_220) begin
                  state <= 8'h4;
                end else begin
                  if (_T_190) begin
                    if (_T_209) begin
                      state <= 8'h3;
                    end else begin
                      state <= _GEN_7;
                    end
                  end else begin
                    state <= _GEN_7;
                  end
                end
              end
            end else begin
              if (_T_220) begin
                state <= 8'h4;
              end else begin
                if (_T_190) begin
                  if (_T_209) begin
                    state <= 8'h3;
                  end else begin
                    state <= _GEN_7;
                  end
                end else begin
                  state <= _GEN_7;
                end
              end
            end
          end
        end else begin
          if (_T_231) begin
            if (_T_256) begin
              state <= 8'h5;
            end else begin
              state <= _GEN_88;
            end
          end else begin
            state <= _GEN_88;
          end
        end
      end
    end
    if (reset) begin
      substate <= 16'h0;
    end else begin
      if (io_en) begin
        if (_T_281) begin
          substate <= _T_204;
        end else begin
          if (_T_231) begin
            if (_T_256) begin
              substate <= 16'h0;
            end else begin
              if (_T_245) begin
                substate <= _T_204;
              end else begin
                if (_T_220) begin
                  substate <= 16'h0;
                end else begin
                  if (_T_190) begin
                    if (_T_209) begin
                      substate <= 16'h0;
                    end else begin
                      if (_T_194) begin
                        substate <= _T_204;
                      end else begin
                        if (_T_186) begin
                          substate <= 16'h0;
                        end else begin
                          if (_T_177) begin
                            substate <= 16'h0;
                          end
                        end
                      end
                    end
                  end else begin
                    if (_T_186) begin
                      substate <= 16'h0;
                    end else begin
                      if (_T_177) begin
                        substate <= 16'h0;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_220) begin
              substate <= 16'h0;
            end else begin
              if (_T_190) begin
                if (_T_209) begin
                  substate <= 16'h0;
                end else begin
                  if (_T_194) begin
                    substate <= _T_204;
                  end else begin
                    if (_T_186) begin
                      substate <= 16'h0;
                    end else begin
                      if (_T_177) begin
                        substate <= 16'h0;
                      end
                    end
                  end
                end
              end else begin
                if (_T_186) begin
                  substate <= 16'h0;
                end else begin
                  if (_T_177) begin
                    substate <= 16'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_en) begin
      if (_T_281) begin
        maxOffsetReg <= _T_315;
      end else begin
        if (_T_231) begin
          if (_T_256) begin
            maxOffsetReg <= 4'h0;
          end
        end
      end
    end
  end
endmodule
