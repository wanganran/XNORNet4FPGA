`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module Memo(
  input         clock,
  input         io_wen,
  input  [7:0]  io_wrAddr,
  input  [17:0] io_wrData,
  input         io_ren,
  input  [7:0]  io_rdAddr,
  output [17:0] io_rdData
);
  reg [17:0] mem [0:255];
  reg [31:0] _GEN_0;
  wire [17:0] mem__T_12_data;
  wire [7:0] mem__T_12_addr;
  wire [17:0] mem__T_10_data;
  wire [7:0] mem__T_10_addr;
  wire  mem__T_10_mask;
  wire  mem__T_10_en;
  reg [7:0] mem__T_12_addr_pipe_0;
  reg [31:0] _GEN_1;
  wire [17:0] _GEN_7;
  assign io_rdData = _GEN_7;
  assign mem__T_12_addr = mem__T_12_addr_pipe_0;
  assign mem__T_12_data = mem[mem__T_12_addr];
  assign mem__T_10_data = io_wrData;
  assign mem__T_10_addr = io_wrAddr;
  assign mem__T_10_mask = io_wen;
  assign mem__T_10_en = io_wen;
  assign _GEN_7 = io_ren ? mem__T_12_data : 18'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    mem[initvar] = _GEN_0[17:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1 = {1{$random}};
  mem__T_12_addr_pipe_0 = _GEN_1[7:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if(mem__T_10_en & mem__T_10_mask) begin
      mem[mem__T_10_addr] <= mem__T_10_data;
    end
    if (io_ren) begin
      mem__T_12_addr_pipe_0 <= io_rdAddr;
    end
  end
endmodule
module AggregateMem(
  input          clock,
  input  [7:0]   io_addr,
  input  [7:0]   io_waddr,
  input  [127:0] io_in,
  output [127:0] io_out,
  input          io_wen,
  input          io_ren
);
  wire  Memo_clock;
  wire  Memo_io_wen;
  wire [7:0] Memo_io_wrAddr;
  wire [17:0] Memo_io_wrData;
  wire  Memo_io_ren;
  wire [7:0] Memo_io_rdAddr;
  wire [17:0] Memo_io_rdData;
  wire  Memo_1_clock;
  wire  Memo_1_io_wen;
  wire [7:0] Memo_1_io_wrAddr;
  wire [17:0] Memo_1_io_wrData;
  wire  Memo_1_io_ren;
  wire [7:0] Memo_1_io_rdAddr;
  wire [17:0] Memo_1_io_rdData;
  wire  Memo_2_clock;
  wire  Memo_2_io_wen;
  wire [7:0] Memo_2_io_wrAddr;
  wire [17:0] Memo_2_io_wrData;
  wire  Memo_2_io_ren;
  wire [7:0] Memo_2_io_rdAddr;
  wire [17:0] Memo_2_io_rdData;
  wire  Memo_3_clock;
  wire  Memo_3_io_wen;
  wire [7:0] Memo_3_io_wrAddr;
  wire [17:0] Memo_3_io_wrData;
  wire  Memo_3_io_ren;
  wire [7:0] Memo_3_io_rdAddr;
  wire [17:0] Memo_3_io_rdData;
  wire  Memo_4_clock;
  wire  Memo_4_io_wen;
  wire [7:0] Memo_4_io_wrAddr;
  wire [17:0] Memo_4_io_wrData;
  wire  Memo_4_io_ren;
  wire [7:0] Memo_4_io_rdAddr;
  wire [17:0] Memo_4_io_rdData;
  wire  Memo_5_clock;
  wire  Memo_5_io_wen;
  wire [7:0] Memo_5_io_wrAddr;
  wire [17:0] Memo_5_io_wrData;
  wire  Memo_5_io_ren;
  wire [7:0] Memo_5_io_rdAddr;
  wire [17:0] Memo_5_io_rdData;
  wire  Memo_6_clock;
  wire  Memo_6_io_wen;
  wire [7:0] Memo_6_io_wrAddr;
  wire [17:0] Memo_6_io_wrData;
  wire  Memo_6_io_ren;
  wire [7:0] Memo_6_io_rdAddr;
  wire [17:0] Memo_6_io_rdData;
  wire  Memo_7_clock;
  wire  Memo_7_io_wen;
  wire [7:0] Memo_7_io_wrAddr;
  wire [17:0] Memo_7_io_wrData;
  wire  Memo_7_io_ren;
  wire [7:0] Memo_7_io_rdAddr;
  wire [17:0] Memo_7_io_rdData;
  wire [15:0] _T_9;
  wire [17:0] _T_10;
  wire [15:0] _T_12;
  wire [17:0] _T_13;
  wire [15:0] _T_15;
  wire [17:0] _T_16;
  wire [15:0] _T_18;
  wire [17:0] _T_19;
  wire [15:0] _T_21;
  wire [17:0] _T_22;
  wire [15:0] _T_24;
  wire [17:0] _T_25;
  wire [15:0] _T_27;
  wire [17:0] _T_28;
  wire [15:0] _T_30;
  wire [17:0] _T_31;
  wire [15:0] _T_32;
  wire [15:0] _T_33;
  wire [15:0] _T_34;
  wire [15:0] _T_35;
  wire [15:0] _T_36;
  wire [15:0] _T_37;
  wire [15:0] _T_38;
  wire [15:0] _T_39;
  wire [31:0] _T_40;
  wire [31:0] _T_41;
  wire [63:0] _T_42;
  wire [31:0] _T_43;
  wire [31:0] _T_44;
  wire [63:0] _T_45;
  wire [127:0] _T_46;
  Memo Memo (
    .clock(Memo_clock),
    .io_wen(Memo_io_wen),
    .io_wrAddr(Memo_io_wrAddr),
    .io_wrData(Memo_io_wrData),
    .io_ren(Memo_io_ren),
    .io_rdAddr(Memo_io_rdAddr),
    .io_rdData(Memo_io_rdData)
  );
  Memo Memo_1 (
    .clock(Memo_1_clock),
    .io_wen(Memo_1_io_wen),
    .io_wrAddr(Memo_1_io_wrAddr),
    .io_wrData(Memo_1_io_wrData),
    .io_ren(Memo_1_io_ren),
    .io_rdAddr(Memo_1_io_rdAddr),
    .io_rdData(Memo_1_io_rdData)
  );
  Memo Memo_2 (
    .clock(Memo_2_clock),
    .io_wen(Memo_2_io_wen),
    .io_wrAddr(Memo_2_io_wrAddr),
    .io_wrData(Memo_2_io_wrData),
    .io_ren(Memo_2_io_ren),
    .io_rdAddr(Memo_2_io_rdAddr),
    .io_rdData(Memo_2_io_rdData)
  );
  Memo Memo_3 (
    .clock(Memo_3_clock),
    .io_wen(Memo_3_io_wen),
    .io_wrAddr(Memo_3_io_wrAddr),
    .io_wrData(Memo_3_io_wrData),
    .io_ren(Memo_3_io_ren),
    .io_rdAddr(Memo_3_io_rdAddr),
    .io_rdData(Memo_3_io_rdData)
  );
  Memo Memo_4 (
    .clock(Memo_4_clock),
    .io_wen(Memo_4_io_wen),
    .io_wrAddr(Memo_4_io_wrAddr),
    .io_wrData(Memo_4_io_wrData),
    .io_ren(Memo_4_io_ren),
    .io_rdAddr(Memo_4_io_rdAddr),
    .io_rdData(Memo_4_io_rdData)
  );
  Memo Memo_5 (
    .clock(Memo_5_clock),
    .io_wen(Memo_5_io_wen),
    .io_wrAddr(Memo_5_io_wrAddr),
    .io_wrData(Memo_5_io_wrData),
    .io_ren(Memo_5_io_ren),
    .io_rdAddr(Memo_5_io_rdAddr),
    .io_rdData(Memo_5_io_rdData)
  );
  Memo Memo_6 (
    .clock(Memo_6_clock),
    .io_wen(Memo_6_io_wen),
    .io_wrAddr(Memo_6_io_wrAddr),
    .io_wrData(Memo_6_io_wrData),
    .io_ren(Memo_6_io_ren),
    .io_rdAddr(Memo_6_io_rdAddr),
    .io_rdData(Memo_6_io_rdData)
  );
  Memo Memo_7 (
    .clock(Memo_7_clock),
    .io_wen(Memo_7_io_wen),
    .io_wrAddr(Memo_7_io_wrAddr),
    .io_wrData(Memo_7_io_wrData),
    .io_ren(Memo_7_io_ren),
    .io_rdAddr(Memo_7_io_rdAddr),
    .io_rdData(Memo_7_io_rdData)
  );
  assign io_out = _T_46;
  assign Memo_clock = clock;
  assign Memo_io_wen = io_wen;
  assign Memo_io_wrAddr = io_waddr;
  assign Memo_io_wrData = _T_10;
  assign Memo_io_ren = io_ren;
  assign Memo_io_rdAddr = io_addr;
  assign Memo_1_clock = clock;
  assign Memo_1_io_wen = io_wen;
  assign Memo_1_io_wrAddr = io_waddr;
  assign Memo_1_io_wrData = _T_13;
  assign Memo_1_io_ren = io_ren;
  assign Memo_1_io_rdAddr = io_addr;
  assign Memo_2_clock = clock;
  assign Memo_2_io_wen = io_wen;
  assign Memo_2_io_wrAddr = io_waddr;
  assign Memo_2_io_wrData = _T_16;
  assign Memo_2_io_ren = io_ren;
  assign Memo_2_io_rdAddr = io_addr;
  assign Memo_3_clock = clock;
  assign Memo_3_io_wen = io_wen;
  assign Memo_3_io_wrAddr = io_waddr;
  assign Memo_3_io_wrData = _T_19;
  assign Memo_3_io_ren = io_ren;
  assign Memo_3_io_rdAddr = io_addr;
  assign Memo_4_clock = clock;
  assign Memo_4_io_wen = io_wen;
  assign Memo_4_io_wrAddr = io_waddr;
  assign Memo_4_io_wrData = _T_22;
  assign Memo_4_io_ren = io_ren;
  assign Memo_4_io_rdAddr = io_addr;
  assign Memo_5_clock = clock;
  assign Memo_5_io_wen = io_wen;
  assign Memo_5_io_wrAddr = io_waddr;
  assign Memo_5_io_wrData = _T_25;
  assign Memo_5_io_ren = io_ren;
  assign Memo_5_io_rdAddr = io_addr;
  assign Memo_6_clock = clock;
  assign Memo_6_io_wen = io_wen;
  assign Memo_6_io_wrAddr = io_waddr;
  assign Memo_6_io_wrData = _T_28;
  assign Memo_6_io_ren = io_ren;
  assign Memo_6_io_rdAddr = io_addr;
  assign Memo_7_clock = clock;
  assign Memo_7_io_wen = io_wen;
  assign Memo_7_io_wrAddr = io_waddr;
  assign Memo_7_io_wrData = _T_31;
  assign Memo_7_io_ren = io_ren;
  assign Memo_7_io_rdAddr = io_addr;
  assign _T_9 = io_in[15:0];
  assign _T_10 = {2'h0,_T_9};
  assign _T_12 = io_in[31:16];
  assign _T_13 = {2'h0,_T_12};
  assign _T_15 = io_in[47:32];
  assign _T_16 = {2'h0,_T_15};
  assign _T_18 = io_in[63:48];
  assign _T_19 = {2'h0,_T_18};
  assign _T_21 = io_in[79:64];
  assign _T_22 = {2'h0,_T_21};
  assign _T_24 = io_in[95:80];
  assign _T_25 = {2'h0,_T_24};
  assign _T_27 = io_in[111:96];
  assign _T_28 = {2'h0,_T_27};
  assign _T_30 = io_in[127:112];
  assign _T_31 = {2'h0,_T_30};
  assign _T_32 = Memo_7_io_rdData[15:0];
  assign _T_33 = Memo_6_io_rdData[15:0];
  assign _T_34 = Memo_5_io_rdData[15:0];
  assign _T_35 = Memo_4_io_rdData[15:0];
  assign _T_36 = Memo_3_io_rdData[15:0];
  assign _T_37 = Memo_2_io_rdData[15:0];
  assign _T_38 = Memo_1_io_rdData[15:0];
  assign _T_39 = Memo_io_rdData[15:0];
  assign _T_40 = {_T_38,_T_39};
  assign _T_41 = {_T_36,_T_37};
  assign _T_42 = {_T_41,_T_40};
  assign _T_43 = {_T_34,_T_35};
  assign _T_44 = {_T_32,_T_33};
  assign _T_45 = {_T_44,_T_43};
  assign _T_46 = {_T_45,_T_42};
endmodule
module BinaryBuffer(
  input          clock,
  input          io_reset,
  input  [3:0]   io_in,
  input  [127:0] io_fastin,
  input          io_push,
  input          io_fastpush,
  output [31:0]  io_out,
  input          io_pop
);
  reg [5:0] wPos;
  reg [31:0] _GEN_2425;
  reg [2:0] rPos;
  reg [31:0] _GEN_2426;
  reg [3:0] mem_0;
  reg [31:0] _GEN_2427;
  reg [3:0] mem_1;
  reg [31:0] _GEN_2428;
  reg [3:0] mem_2;
  reg [31:0] _GEN_2429;
  reg [3:0] mem_3;
  reg [31:0] _GEN_2430;
  reg [3:0] mem_4;
  reg [31:0] _GEN_2431;
  reg [3:0] mem_5;
  reg [31:0] _GEN_2432;
  reg [3:0] mem_6;
  reg [31:0] _GEN_2433;
  reg [3:0] mem_7;
  reg [31:0] _GEN_2434;
  reg [3:0] mem_8;
  reg [31:0] _GEN_2435;
  reg [3:0] mem_9;
  reg [31:0] _GEN_2436;
  reg [3:0] mem_10;
  reg [31:0] _GEN_2437;
  reg [3:0] mem_11;
  reg [31:0] _GEN_2438;
  reg [3:0] mem_12;
  reg [31:0] _GEN_2439;
  reg [3:0] mem_13;
  reg [31:0] _GEN_2440;
  reg [3:0] mem_14;
  reg [31:0] _GEN_2441;
  reg [3:0] mem_15;
  reg [31:0] _GEN_2442;
  reg [3:0] mem_16;
  reg [31:0] _GEN_2443;
  reg [3:0] mem_17;
  reg [31:0] _GEN_2444;
  reg [3:0] mem_18;
  reg [31:0] _GEN_2445;
  reg [3:0] mem_19;
  reg [31:0] _GEN_2446;
  reg [3:0] mem_20;
  reg [31:0] _GEN_2447;
  reg [3:0] mem_21;
  reg [31:0] _GEN_2448;
  reg [3:0] mem_22;
  reg [31:0] _GEN_2449;
  reg [3:0] mem_23;
  reg [31:0] _GEN_2450;
  reg [3:0] mem_24;
  reg [31:0] _GEN_2451;
  reg [3:0] mem_25;
  reg [31:0] _GEN_2452;
  reg [3:0] mem_26;
  reg [31:0] _GEN_2453;
  reg [3:0] mem_27;
  reg [31:0] _GEN_2454;
  reg [3:0] mem_28;
  reg [31:0] _GEN_2455;
  reg [3:0] mem_29;
  reg [31:0] _GEN_2456;
  reg [3:0] mem_30;
  reg [31:0] _GEN_2457;
  reg [3:0] mem_31;
  reg [31:0] _GEN_2458;
  reg [3:0] mem_32;
  reg [31:0] _GEN_2459;
  reg [3:0] mem_33;
  reg [31:0] _GEN_2460;
  reg [3:0] mem_34;
  reg [31:0] _GEN_2461;
  reg [3:0] mem_35;
  reg [31:0] _GEN_2462;
  reg [3:0] mem_36;
  reg [31:0] _GEN_2463;
  reg [3:0] mem_37;
  reg [31:0] _GEN_2464;
  reg [3:0] mem_38;
  reg [31:0] _GEN_2465;
  reg [3:0] mem_39;
  reg [31:0] _GEN_2466;
  reg [3:0] mem_40;
  reg [31:0] _GEN_2467;
  reg [3:0] mem_41;
  reg [31:0] _GEN_2468;
  reg [3:0] mem_42;
  reg [31:0] _GEN_2469;
  reg [3:0] mem_43;
  reg [31:0] _GEN_2470;
  reg [3:0] mem_44;
  reg [31:0] _GEN_2471;
  reg [3:0] mem_45;
  reg [31:0] _GEN_2472;
  reg [3:0] mem_46;
  reg [31:0] _GEN_2473;
  reg [3:0] mem_47;
  reg [31:0] _GEN_2474;
  reg [3:0] mem_48;
  reg [31:0] _GEN_2475;
  reg [3:0] mem_49;
  reg [31:0] _GEN_2476;
  reg [3:0] mem_50;
  reg [31:0] _GEN_2477;
  reg [3:0] mem_51;
  reg [31:0] _GEN_2478;
  reg [3:0] mem_52;
  reg [31:0] _GEN_2479;
  reg [3:0] mem_53;
  reg [31:0] _GEN_2480;
  reg [3:0] mem_54;
  reg [31:0] _GEN_2481;
  reg [3:0] mem_55;
  reg [31:0] _GEN_2482;
  reg [3:0] mem_56;
  reg [31:0] _GEN_2483;
  reg [3:0] mem_57;
  reg [31:0] _GEN_2484;
  reg [3:0] mem_58;
  reg [31:0] _GEN_2485;
  reg [3:0] mem_59;
  reg [31:0] _GEN_2486;
  reg [3:0] mem_60;
  reg [31:0] _GEN_2487;
  reg [3:0] mem_61;
  reg [31:0] _GEN_2488;
  reg [3:0] mem_62;
  reg [31:0] _GEN_2489;
  reg [3:0] mem_63;
  reg [31:0] _GEN_2490;
  wire [7:0] _T_80;
  wire [7:0] _T_81;
  wire [15:0] _T_82;
  wire [7:0] _T_83;
  wire [7:0] _T_84;
  wire [15:0] _T_85;
  wire [31:0] _T_86;
  wire [7:0] _T_87;
  wire [7:0] _T_88;
  wire [15:0] _T_89;
  wire [7:0] _T_90;
  wire [7:0] _T_91;
  wire [15:0] _T_92;
  wire [31:0] _T_93;
  wire [7:0] _T_94;
  wire [7:0] _T_95;
  wire [15:0] _T_96;
  wire [7:0] _T_97;
  wire [7:0] _T_98;
  wire [15:0] _T_99;
  wire [31:0] _T_100;
  wire [7:0] _T_101;
  wire [7:0] _T_102;
  wire [15:0] _T_103;
  wire [7:0] _T_104;
  wire [7:0] _T_105;
  wire [15:0] _T_106;
  wire [31:0] _T_107;
  wire [7:0] _T_108;
  wire [7:0] _T_109;
  wire [15:0] _T_110;
  wire [7:0] _T_111;
  wire [7:0] _T_112;
  wire [15:0] _T_113;
  wire [31:0] _T_114;
  wire [7:0] _T_115;
  wire [7:0] _T_116;
  wire [15:0] _T_117;
  wire [7:0] _T_118;
  wire [7:0] _T_119;
  wire [15:0] _T_120;
  wire [31:0] _T_121;
  wire [7:0] _T_122;
  wire [7:0] _T_123;
  wire [15:0] _T_124;
  wire [7:0] _T_125;
  wire [7:0] _T_126;
  wire [15:0] _T_127;
  wire [31:0] _T_128;
  wire [7:0] _T_129;
  wire [7:0] _T_130;
  wire [15:0] _T_131;
  wire [7:0] _T_132;
  wire [7:0] _T_133;
  wire [15:0] _T_134;
  wire [31:0] _T_135;
  wire [31:0] catMem_0;
  wire [31:0] catMem_1;
  wire [31:0] catMem_2;
  wire [31:0] catMem_3;
  wire [31:0] catMem_4;
  wire [31:0] catMem_5;
  wire [31:0] catMem_6;
  wire [31:0] catMem_7;
  wire  _T_149;
  wire  _T_150;
  wire [6:0] _T_152;
  wire [5:0] _T_153;
  wire [3:0] _T_155;
  wire [3:0] _GEN_0;
  wire [3:0] _GEN_34;
  wire [3:0] _GEN_35;
  wire [3:0] _GEN_36;
  wire [3:0] _GEN_37;
  wire [3:0] _GEN_38;
  wire [3:0] _GEN_39;
  wire [3:0] _GEN_40;
  wire [3:0] _GEN_41;
  wire [3:0] _GEN_42;
  wire [3:0] _GEN_43;
  wire [3:0] _GEN_44;
  wire [3:0] _GEN_45;
  wire [3:0] _GEN_46;
  wire [3:0] _GEN_47;
  wire [3:0] _GEN_48;
  wire [3:0] _GEN_49;
  wire [3:0] _GEN_50;
  wire [3:0] _GEN_51;
  wire [3:0] _GEN_52;
  wire [3:0] _GEN_53;
  wire [3:0] _GEN_54;
  wire [3:0] _GEN_55;
  wire [3:0] _GEN_56;
  wire [3:0] _GEN_57;
  wire [3:0] _GEN_58;
  wire [3:0] _GEN_59;
  wire [3:0] _GEN_60;
  wire [3:0] _GEN_61;
  wire [3:0] _GEN_62;
  wire [3:0] _GEN_63;
  wire [3:0] _GEN_64;
  wire [3:0] _GEN_65;
  wire [3:0] _GEN_66;
  wire [3:0] _GEN_67;
  wire [3:0] _GEN_68;
  wire [3:0] _GEN_69;
  wire [3:0] _GEN_70;
  wire [3:0] _GEN_71;
  wire [3:0] _GEN_72;
  wire [3:0] _GEN_73;
  wire [3:0] _GEN_74;
  wire [3:0] _GEN_75;
  wire [3:0] _GEN_76;
  wire [3:0] _GEN_77;
  wire [3:0] _GEN_78;
  wire [3:0] _GEN_79;
  wire [3:0] _GEN_80;
  wire [3:0] _GEN_81;
  wire [3:0] _GEN_82;
  wire [3:0] _GEN_83;
  wire [3:0] _GEN_84;
  wire [3:0] _GEN_85;
  wire [3:0] _GEN_86;
  wire [3:0] _GEN_87;
  wire [3:0] _GEN_88;
  wire [3:0] _GEN_89;
  wire [3:0] _GEN_90;
  wire [3:0] _GEN_91;
  wire [3:0] _GEN_92;
  wire [3:0] _GEN_93;
  wire [3:0] _GEN_94;
  wire [3:0] _GEN_95;
  wire [3:0] _GEN_96;
  wire [3:0] _GEN_97;
  wire [6:0] _T_157;
  wire [5:0] _T_158;
  wire [3:0] _T_160;
  wire [3:0] _GEN_1;
  wire [3:0] _GEN_98;
  wire [3:0] _GEN_99;
  wire [3:0] _GEN_100;
  wire [3:0] _GEN_101;
  wire [3:0] _GEN_102;
  wire [3:0] _GEN_103;
  wire [3:0] _GEN_104;
  wire [3:0] _GEN_105;
  wire [3:0] _GEN_106;
  wire [3:0] _GEN_107;
  wire [3:0] _GEN_108;
  wire [3:0] _GEN_109;
  wire [3:0] _GEN_110;
  wire [3:0] _GEN_111;
  wire [3:0] _GEN_112;
  wire [3:0] _GEN_113;
  wire [3:0] _GEN_114;
  wire [3:0] _GEN_115;
  wire [3:0] _GEN_116;
  wire [3:0] _GEN_117;
  wire [3:0] _GEN_118;
  wire [3:0] _GEN_119;
  wire [3:0] _GEN_120;
  wire [3:0] _GEN_121;
  wire [3:0] _GEN_122;
  wire [3:0] _GEN_123;
  wire [3:0] _GEN_124;
  wire [3:0] _GEN_125;
  wire [3:0] _GEN_126;
  wire [3:0] _GEN_127;
  wire [3:0] _GEN_128;
  wire [3:0] _GEN_129;
  wire [3:0] _GEN_130;
  wire [3:0] _GEN_131;
  wire [3:0] _GEN_132;
  wire [3:0] _GEN_133;
  wire [3:0] _GEN_134;
  wire [3:0] _GEN_135;
  wire [3:0] _GEN_136;
  wire [3:0] _GEN_137;
  wire [3:0] _GEN_138;
  wire [3:0] _GEN_139;
  wire [3:0] _GEN_140;
  wire [3:0] _GEN_141;
  wire [3:0] _GEN_142;
  wire [3:0] _GEN_143;
  wire [3:0] _GEN_144;
  wire [3:0] _GEN_145;
  wire [3:0] _GEN_146;
  wire [3:0] _GEN_147;
  wire [3:0] _GEN_148;
  wire [3:0] _GEN_149;
  wire [3:0] _GEN_150;
  wire [3:0] _GEN_151;
  wire [3:0] _GEN_152;
  wire [3:0] _GEN_153;
  wire [3:0] _GEN_154;
  wire [3:0] _GEN_155;
  wire [3:0] _GEN_156;
  wire [3:0] _GEN_157;
  wire [3:0] _GEN_158;
  wire [3:0] _GEN_159;
  wire [3:0] _GEN_160;
  wire [3:0] _GEN_161;
  wire [6:0] _T_162;
  wire [5:0] _T_163;
  wire [3:0] _T_165;
  wire [3:0] _GEN_2;
  wire [3:0] _GEN_162;
  wire [3:0] _GEN_163;
  wire [3:0] _GEN_164;
  wire [3:0] _GEN_165;
  wire [3:0] _GEN_166;
  wire [3:0] _GEN_167;
  wire [3:0] _GEN_168;
  wire [3:0] _GEN_169;
  wire [3:0] _GEN_170;
  wire [3:0] _GEN_171;
  wire [3:0] _GEN_172;
  wire [3:0] _GEN_173;
  wire [3:0] _GEN_174;
  wire [3:0] _GEN_175;
  wire [3:0] _GEN_176;
  wire [3:0] _GEN_177;
  wire [3:0] _GEN_178;
  wire [3:0] _GEN_179;
  wire [3:0] _GEN_180;
  wire [3:0] _GEN_181;
  wire [3:0] _GEN_182;
  wire [3:0] _GEN_183;
  wire [3:0] _GEN_184;
  wire [3:0] _GEN_185;
  wire [3:0] _GEN_186;
  wire [3:0] _GEN_187;
  wire [3:0] _GEN_188;
  wire [3:0] _GEN_189;
  wire [3:0] _GEN_190;
  wire [3:0] _GEN_191;
  wire [3:0] _GEN_192;
  wire [3:0] _GEN_193;
  wire [3:0] _GEN_194;
  wire [3:0] _GEN_195;
  wire [3:0] _GEN_196;
  wire [3:0] _GEN_197;
  wire [3:0] _GEN_198;
  wire [3:0] _GEN_199;
  wire [3:0] _GEN_200;
  wire [3:0] _GEN_201;
  wire [3:0] _GEN_202;
  wire [3:0] _GEN_203;
  wire [3:0] _GEN_204;
  wire [3:0] _GEN_205;
  wire [3:0] _GEN_206;
  wire [3:0] _GEN_207;
  wire [3:0] _GEN_208;
  wire [3:0] _GEN_209;
  wire [3:0] _GEN_210;
  wire [3:0] _GEN_211;
  wire [3:0] _GEN_212;
  wire [3:0] _GEN_213;
  wire [3:0] _GEN_214;
  wire [3:0] _GEN_215;
  wire [3:0] _GEN_216;
  wire [3:0] _GEN_217;
  wire [3:0] _GEN_218;
  wire [3:0] _GEN_219;
  wire [3:0] _GEN_220;
  wire [3:0] _GEN_221;
  wire [3:0] _GEN_222;
  wire [3:0] _GEN_223;
  wire [3:0] _GEN_224;
  wire [3:0] _GEN_225;
  wire [6:0] _T_167;
  wire [5:0] _T_168;
  wire [3:0] _T_170;
  wire [3:0] _GEN_3;
  wire [3:0] _GEN_226;
  wire [3:0] _GEN_227;
  wire [3:0] _GEN_228;
  wire [3:0] _GEN_229;
  wire [3:0] _GEN_230;
  wire [3:0] _GEN_231;
  wire [3:0] _GEN_232;
  wire [3:0] _GEN_233;
  wire [3:0] _GEN_234;
  wire [3:0] _GEN_235;
  wire [3:0] _GEN_236;
  wire [3:0] _GEN_237;
  wire [3:0] _GEN_238;
  wire [3:0] _GEN_239;
  wire [3:0] _GEN_240;
  wire [3:0] _GEN_241;
  wire [3:0] _GEN_242;
  wire [3:0] _GEN_243;
  wire [3:0] _GEN_244;
  wire [3:0] _GEN_245;
  wire [3:0] _GEN_246;
  wire [3:0] _GEN_247;
  wire [3:0] _GEN_248;
  wire [3:0] _GEN_249;
  wire [3:0] _GEN_250;
  wire [3:0] _GEN_251;
  wire [3:0] _GEN_252;
  wire [3:0] _GEN_253;
  wire [3:0] _GEN_254;
  wire [3:0] _GEN_255;
  wire [3:0] _GEN_256;
  wire [3:0] _GEN_257;
  wire [3:0] _GEN_258;
  wire [3:0] _GEN_259;
  wire [3:0] _GEN_260;
  wire [3:0] _GEN_261;
  wire [3:0] _GEN_262;
  wire [3:0] _GEN_263;
  wire [3:0] _GEN_264;
  wire [3:0] _GEN_265;
  wire [3:0] _GEN_266;
  wire [3:0] _GEN_267;
  wire [3:0] _GEN_268;
  wire [3:0] _GEN_269;
  wire [3:0] _GEN_270;
  wire [3:0] _GEN_271;
  wire [3:0] _GEN_272;
  wire [3:0] _GEN_273;
  wire [3:0] _GEN_274;
  wire [3:0] _GEN_275;
  wire [3:0] _GEN_276;
  wire [3:0] _GEN_277;
  wire [3:0] _GEN_278;
  wire [3:0] _GEN_279;
  wire [3:0] _GEN_280;
  wire [3:0] _GEN_281;
  wire [3:0] _GEN_282;
  wire [3:0] _GEN_283;
  wire [3:0] _GEN_284;
  wire [3:0] _GEN_285;
  wire [3:0] _GEN_286;
  wire [3:0] _GEN_287;
  wire [3:0] _GEN_288;
  wire [3:0] _GEN_289;
  wire [6:0] _T_172;
  wire [5:0] _T_173;
  wire [3:0] _T_175;
  wire [3:0] _GEN_4;
  wire [3:0] _GEN_290;
  wire [3:0] _GEN_291;
  wire [3:0] _GEN_292;
  wire [3:0] _GEN_293;
  wire [3:0] _GEN_294;
  wire [3:0] _GEN_295;
  wire [3:0] _GEN_296;
  wire [3:0] _GEN_297;
  wire [3:0] _GEN_298;
  wire [3:0] _GEN_299;
  wire [3:0] _GEN_300;
  wire [3:0] _GEN_301;
  wire [3:0] _GEN_302;
  wire [3:0] _GEN_303;
  wire [3:0] _GEN_304;
  wire [3:0] _GEN_305;
  wire [3:0] _GEN_306;
  wire [3:0] _GEN_307;
  wire [3:0] _GEN_308;
  wire [3:0] _GEN_309;
  wire [3:0] _GEN_310;
  wire [3:0] _GEN_311;
  wire [3:0] _GEN_312;
  wire [3:0] _GEN_313;
  wire [3:0] _GEN_314;
  wire [3:0] _GEN_315;
  wire [3:0] _GEN_316;
  wire [3:0] _GEN_317;
  wire [3:0] _GEN_318;
  wire [3:0] _GEN_319;
  wire [3:0] _GEN_320;
  wire [3:0] _GEN_321;
  wire [3:0] _GEN_322;
  wire [3:0] _GEN_323;
  wire [3:0] _GEN_324;
  wire [3:0] _GEN_325;
  wire [3:0] _GEN_326;
  wire [3:0] _GEN_327;
  wire [3:0] _GEN_328;
  wire [3:0] _GEN_329;
  wire [3:0] _GEN_330;
  wire [3:0] _GEN_331;
  wire [3:0] _GEN_332;
  wire [3:0] _GEN_333;
  wire [3:0] _GEN_334;
  wire [3:0] _GEN_335;
  wire [3:0] _GEN_336;
  wire [3:0] _GEN_337;
  wire [3:0] _GEN_338;
  wire [3:0] _GEN_339;
  wire [3:0] _GEN_340;
  wire [3:0] _GEN_341;
  wire [3:0] _GEN_342;
  wire [3:0] _GEN_343;
  wire [3:0] _GEN_344;
  wire [3:0] _GEN_345;
  wire [3:0] _GEN_346;
  wire [3:0] _GEN_347;
  wire [3:0] _GEN_348;
  wire [3:0] _GEN_349;
  wire [3:0] _GEN_350;
  wire [3:0] _GEN_351;
  wire [3:0] _GEN_352;
  wire [3:0] _GEN_353;
  wire [6:0] _T_177;
  wire [5:0] _T_178;
  wire [3:0] _T_180;
  wire [3:0] _GEN_5;
  wire [3:0] _GEN_354;
  wire [3:0] _GEN_355;
  wire [3:0] _GEN_356;
  wire [3:0] _GEN_357;
  wire [3:0] _GEN_358;
  wire [3:0] _GEN_359;
  wire [3:0] _GEN_360;
  wire [3:0] _GEN_361;
  wire [3:0] _GEN_362;
  wire [3:0] _GEN_363;
  wire [3:0] _GEN_364;
  wire [3:0] _GEN_365;
  wire [3:0] _GEN_366;
  wire [3:0] _GEN_367;
  wire [3:0] _GEN_368;
  wire [3:0] _GEN_369;
  wire [3:0] _GEN_370;
  wire [3:0] _GEN_371;
  wire [3:0] _GEN_372;
  wire [3:0] _GEN_373;
  wire [3:0] _GEN_374;
  wire [3:0] _GEN_375;
  wire [3:0] _GEN_376;
  wire [3:0] _GEN_377;
  wire [3:0] _GEN_378;
  wire [3:0] _GEN_379;
  wire [3:0] _GEN_380;
  wire [3:0] _GEN_381;
  wire [3:0] _GEN_382;
  wire [3:0] _GEN_383;
  wire [3:0] _GEN_384;
  wire [3:0] _GEN_385;
  wire [3:0] _GEN_386;
  wire [3:0] _GEN_387;
  wire [3:0] _GEN_388;
  wire [3:0] _GEN_389;
  wire [3:0] _GEN_390;
  wire [3:0] _GEN_391;
  wire [3:0] _GEN_392;
  wire [3:0] _GEN_393;
  wire [3:0] _GEN_394;
  wire [3:0] _GEN_395;
  wire [3:0] _GEN_396;
  wire [3:0] _GEN_397;
  wire [3:0] _GEN_398;
  wire [3:0] _GEN_399;
  wire [3:0] _GEN_400;
  wire [3:0] _GEN_401;
  wire [3:0] _GEN_402;
  wire [3:0] _GEN_403;
  wire [3:0] _GEN_404;
  wire [3:0] _GEN_405;
  wire [3:0] _GEN_406;
  wire [3:0] _GEN_407;
  wire [3:0] _GEN_408;
  wire [3:0] _GEN_409;
  wire [3:0] _GEN_410;
  wire [3:0] _GEN_411;
  wire [3:0] _GEN_412;
  wire [3:0] _GEN_413;
  wire [3:0] _GEN_414;
  wire [3:0] _GEN_415;
  wire [3:0] _GEN_416;
  wire [3:0] _GEN_417;
  wire [6:0] _T_182;
  wire [5:0] _T_183;
  wire [3:0] _T_185;
  wire [3:0] _GEN_6;
  wire [3:0] _GEN_418;
  wire [3:0] _GEN_419;
  wire [3:0] _GEN_420;
  wire [3:0] _GEN_421;
  wire [3:0] _GEN_422;
  wire [3:0] _GEN_423;
  wire [3:0] _GEN_424;
  wire [3:0] _GEN_425;
  wire [3:0] _GEN_426;
  wire [3:0] _GEN_427;
  wire [3:0] _GEN_428;
  wire [3:0] _GEN_429;
  wire [3:0] _GEN_430;
  wire [3:0] _GEN_431;
  wire [3:0] _GEN_432;
  wire [3:0] _GEN_433;
  wire [3:0] _GEN_434;
  wire [3:0] _GEN_435;
  wire [3:0] _GEN_436;
  wire [3:0] _GEN_437;
  wire [3:0] _GEN_438;
  wire [3:0] _GEN_439;
  wire [3:0] _GEN_440;
  wire [3:0] _GEN_441;
  wire [3:0] _GEN_442;
  wire [3:0] _GEN_443;
  wire [3:0] _GEN_444;
  wire [3:0] _GEN_445;
  wire [3:0] _GEN_446;
  wire [3:0] _GEN_447;
  wire [3:0] _GEN_448;
  wire [3:0] _GEN_449;
  wire [3:0] _GEN_450;
  wire [3:0] _GEN_451;
  wire [3:0] _GEN_452;
  wire [3:0] _GEN_453;
  wire [3:0] _GEN_454;
  wire [3:0] _GEN_455;
  wire [3:0] _GEN_456;
  wire [3:0] _GEN_457;
  wire [3:0] _GEN_458;
  wire [3:0] _GEN_459;
  wire [3:0] _GEN_460;
  wire [3:0] _GEN_461;
  wire [3:0] _GEN_462;
  wire [3:0] _GEN_463;
  wire [3:0] _GEN_464;
  wire [3:0] _GEN_465;
  wire [3:0] _GEN_466;
  wire [3:0] _GEN_467;
  wire [3:0] _GEN_468;
  wire [3:0] _GEN_469;
  wire [3:0] _GEN_470;
  wire [3:0] _GEN_471;
  wire [3:0] _GEN_472;
  wire [3:0] _GEN_473;
  wire [3:0] _GEN_474;
  wire [3:0] _GEN_475;
  wire [3:0] _GEN_476;
  wire [3:0] _GEN_477;
  wire [3:0] _GEN_478;
  wire [3:0] _GEN_479;
  wire [3:0] _GEN_480;
  wire [3:0] _GEN_481;
  wire [6:0] _T_187;
  wire [5:0] _T_188;
  wire [3:0] _T_190;
  wire [3:0] _GEN_7;
  wire [3:0] _GEN_482;
  wire [3:0] _GEN_483;
  wire [3:0] _GEN_484;
  wire [3:0] _GEN_485;
  wire [3:0] _GEN_486;
  wire [3:0] _GEN_487;
  wire [3:0] _GEN_488;
  wire [3:0] _GEN_489;
  wire [3:0] _GEN_490;
  wire [3:0] _GEN_491;
  wire [3:0] _GEN_492;
  wire [3:0] _GEN_493;
  wire [3:0] _GEN_494;
  wire [3:0] _GEN_495;
  wire [3:0] _GEN_496;
  wire [3:0] _GEN_497;
  wire [3:0] _GEN_498;
  wire [3:0] _GEN_499;
  wire [3:0] _GEN_500;
  wire [3:0] _GEN_501;
  wire [3:0] _GEN_502;
  wire [3:0] _GEN_503;
  wire [3:0] _GEN_504;
  wire [3:0] _GEN_505;
  wire [3:0] _GEN_506;
  wire [3:0] _GEN_507;
  wire [3:0] _GEN_508;
  wire [3:0] _GEN_509;
  wire [3:0] _GEN_510;
  wire [3:0] _GEN_511;
  wire [3:0] _GEN_512;
  wire [3:0] _GEN_513;
  wire [3:0] _GEN_514;
  wire [3:0] _GEN_515;
  wire [3:0] _GEN_516;
  wire [3:0] _GEN_517;
  wire [3:0] _GEN_518;
  wire [3:0] _GEN_519;
  wire [3:0] _GEN_520;
  wire [3:0] _GEN_521;
  wire [3:0] _GEN_522;
  wire [3:0] _GEN_523;
  wire [3:0] _GEN_524;
  wire [3:0] _GEN_525;
  wire [3:0] _GEN_526;
  wire [3:0] _GEN_527;
  wire [3:0] _GEN_528;
  wire [3:0] _GEN_529;
  wire [3:0] _GEN_530;
  wire [3:0] _GEN_531;
  wire [3:0] _GEN_532;
  wire [3:0] _GEN_533;
  wire [3:0] _GEN_534;
  wire [3:0] _GEN_535;
  wire [3:0] _GEN_536;
  wire [3:0] _GEN_537;
  wire [3:0] _GEN_538;
  wire [3:0] _GEN_539;
  wire [3:0] _GEN_540;
  wire [3:0] _GEN_541;
  wire [3:0] _GEN_542;
  wire [3:0] _GEN_543;
  wire [3:0] _GEN_544;
  wire [3:0] _GEN_545;
  wire [6:0] _T_192;
  wire [5:0] _T_193;
  wire [3:0] _T_195;
  wire [3:0] _GEN_8;
  wire [3:0] _GEN_546;
  wire [3:0] _GEN_547;
  wire [3:0] _GEN_548;
  wire [3:0] _GEN_549;
  wire [3:0] _GEN_550;
  wire [3:0] _GEN_551;
  wire [3:0] _GEN_552;
  wire [3:0] _GEN_553;
  wire [3:0] _GEN_554;
  wire [3:0] _GEN_555;
  wire [3:0] _GEN_556;
  wire [3:0] _GEN_557;
  wire [3:0] _GEN_558;
  wire [3:0] _GEN_559;
  wire [3:0] _GEN_560;
  wire [3:0] _GEN_561;
  wire [3:0] _GEN_562;
  wire [3:0] _GEN_563;
  wire [3:0] _GEN_564;
  wire [3:0] _GEN_565;
  wire [3:0] _GEN_566;
  wire [3:0] _GEN_567;
  wire [3:0] _GEN_568;
  wire [3:0] _GEN_569;
  wire [3:0] _GEN_570;
  wire [3:0] _GEN_571;
  wire [3:0] _GEN_572;
  wire [3:0] _GEN_573;
  wire [3:0] _GEN_574;
  wire [3:0] _GEN_575;
  wire [3:0] _GEN_576;
  wire [3:0] _GEN_577;
  wire [3:0] _GEN_578;
  wire [3:0] _GEN_579;
  wire [3:0] _GEN_580;
  wire [3:0] _GEN_581;
  wire [3:0] _GEN_582;
  wire [3:0] _GEN_583;
  wire [3:0] _GEN_584;
  wire [3:0] _GEN_585;
  wire [3:0] _GEN_586;
  wire [3:0] _GEN_587;
  wire [3:0] _GEN_588;
  wire [3:0] _GEN_589;
  wire [3:0] _GEN_590;
  wire [3:0] _GEN_591;
  wire [3:0] _GEN_592;
  wire [3:0] _GEN_593;
  wire [3:0] _GEN_594;
  wire [3:0] _GEN_595;
  wire [3:0] _GEN_596;
  wire [3:0] _GEN_597;
  wire [3:0] _GEN_598;
  wire [3:0] _GEN_599;
  wire [3:0] _GEN_600;
  wire [3:0] _GEN_601;
  wire [3:0] _GEN_602;
  wire [3:0] _GEN_603;
  wire [3:0] _GEN_604;
  wire [3:0] _GEN_605;
  wire [3:0] _GEN_606;
  wire [3:0] _GEN_607;
  wire [3:0] _GEN_608;
  wire [3:0] _GEN_609;
  wire [6:0] _T_197;
  wire [5:0] _T_198;
  wire [3:0] _T_200;
  wire [3:0] _GEN_9;
  wire [3:0] _GEN_610;
  wire [3:0] _GEN_611;
  wire [3:0] _GEN_612;
  wire [3:0] _GEN_613;
  wire [3:0] _GEN_614;
  wire [3:0] _GEN_615;
  wire [3:0] _GEN_616;
  wire [3:0] _GEN_617;
  wire [3:0] _GEN_618;
  wire [3:0] _GEN_619;
  wire [3:0] _GEN_620;
  wire [3:0] _GEN_621;
  wire [3:0] _GEN_622;
  wire [3:0] _GEN_623;
  wire [3:0] _GEN_624;
  wire [3:0] _GEN_625;
  wire [3:0] _GEN_626;
  wire [3:0] _GEN_627;
  wire [3:0] _GEN_628;
  wire [3:0] _GEN_629;
  wire [3:0] _GEN_630;
  wire [3:0] _GEN_631;
  wire [3:0] _GEN_632;
  wire [3:0] _GEN_633;
  wire [3:0] _GEN_634;
  wire [3:0] _GEN_635;
  wire [3:0] _GEN_636;
  wire [3:0] _GEN_637;
  wire [3:0] _GEN_638;
  wire [3:0] _GEN_639;
  wire [3:0] _GEN_640;
  wire [3:0] _GEN_641;
  wire [3:0] _GEN_642;
  wire [3:0] _GEN_643;
  wire [3:0] _GEN_644;
  wire [3:0] _GEN_645;
  wire [3:0] _GEN_646;
  wire [3:0] _GEN_647;
  wire [3:0] _GEN_648;
  wire [3:0] _GEN_649;
  wire [3:0] _GEN_650;
  wire [3:0] _GEN_651;
  wire [3:0] _GEN_652;
  wire [3:0] _GEN_653;
  wire [3:0] _GEN_654;
  wire [3:0] _GEN_655;
  wire [3:0] _GEN_656;
  wire [3:0] _GEN_657;
  wire [3:0] _GEN_658;
  wire [3:0] _GEN_659;
  wire [3:0] _GEN_660;
  wire [3:0] _GEN_661;
  wire [3:0] _GEN_662;
  wire [3:0] _GEN_663;
  wire [3:0] _GEN_664;
  wire [3:0] _GEN_665;
  wire [3:0] _GEN_666;
  wire [3:0] _GEN_667;
  wire [3:0] _GEN_668;
  wire [3:0] _GEN_669;
  wire [3:0] _GEN_670;
  wire [3:0] _GEN_671;
  wire [3:0] _GEN_672;
  wire [3:0] _GEN_673;
  wire [6:0] _T_202;
  wire [5:0] _T_203;
  wire [3:0] _T_205;
  wire [3:0] _GEN_10;
  wire [3:0] _GEN_674;
  wire [3:0] _GEN_675;
  wire [3:0] _GEN_676;
  wire [3:0] _GEN_677;
  wire [3:0] _GEN_678;
  wire [3:0] _GEN_679;
  wire [3:0] _GEN_680;
  wire [3:0] _GEN_681;
  wire [3:0] _GEN_682;
  wire [3:0] _GEN_683;
  wire [3:0] _GEN_684;
  wire [3:0] _GEN_685;
  wire [3:0] _GEN_686;
  wire [3:0] _GEN_687;
  wire [3:0] _GEN_688;
  wire [3:0] _GEN_689;
  wire [3:0] _GEN_690;
  wire [3:0] _GEN_691;
  wire [3:0] _GEN_692;
  wire [3:0] _GEN_693;
  wire [3:0] _GEN_694;
  wire [3:0] _GEN_695;
  wire [3:0] _GEN_696;
  wire [3:0] _GEN_697;
  wire [3:0] _GEN_698;
  wire [3:0] _GEN_699;
  wire [3:0] _GEN_700;
  wire [3:0] _GEN_701;
  wire [3:0] _GEN_702;
  wire [3:0] _GEN_703;
  wire [3:0] _GEN_704;
  wire [3:0] _GEN_705;
  wire [3:0] _GEN_706;
  wire [3:0] _GEN_707;
  wire [3:0] _GEN_708;
  wire [3:0] _GEN_709;
  wire [3:0] _GEN_710;
  wire [3:0] _GEN_711;
  wire [3:0] _GEN_712;
  wire [3:0] _GEN_713;
  wire [3:0] _GEN_714;
  wire [3:0] _GEN_715;
  wire [3:0] _GEN_716;
  wire [3:0] _GEN_717;
  wire [3:0] _GEN_718;
  wire [3:0] _GEN_719;
  wire [3:0] _GEN_720;
  wire [3:0] _GEN_721;
  wire [3:0] _GEN_722;
  wire [3:0] _GEN_723;
  wire [3:0] _GEN_724;
  wire [3:0] _GEN_725;
  wire [3:0] _GEN_726;
  wire [3:0] _GEN_727;
  wire [3:0] _GEN_728;
  wire [3:0] _GEN_729;
  wire [3:0] _GEN_730;
  wire [3:0] _GEN_731;
  wire [3:0] _GEN_732;
  wire [3:0] _GEN_733;
  wire [3:0] _GEN_734;
  wire [3:0] _GEN_735;
  wire [3:0] _GEN_736;
  wire [3:0] _GEN_737;
  wire [6:0] _T_207;
  wire [5:0] _T_208;
  wire [3:0] _T_210;
  wire [3:0] _GEN_11;
  wire [3:0] _GEN_738;
  wire [3:0] _GEN_739;
  wire [3:0] _GEN_740;
  wire [3:0] _GEN_741;
  wire [3:0] _GEN_742;
  wire [3:0] _GEN_743;
  wire [3:0] _GEN_744;
  wire [3:0] _GEN_745;
  wire [3:0] _GEN_746;
  wire [3:0] _GEN_747;
  wire [3:0] _GEN_748;
  wire [3:0] _GEN_749;
  wire [3:0] _GEN_750;
  wire [3:0] _GEN_751;
  wire [3:0] _GEN_752;
  wire [3:0] _GEN_753;
  wire [3:0] _GEN_754;
  wire [3:0] _GEN_755;
  wire [3:0] _GEN_756;
  wire [3:0] _GEN_757;
  wire [3:0] _GEN_758;
  wire [3:0] _GEN_759;
  wire [3:0] _GEN_760;
  wire [3:0] _GEN_761;
  wire [3:0] _GEN_762;
  wire [3:0] _GEN_763;
  wire [3:0] _GEN_764;
  wire [3:0] _GEN_765;
  wire [3:0] _GEN_766;
  wire [3:0] _GEN_767;
  wire [3:0] _GEN_768;
  wire [3:0] _GEN_769;
  wire [3:0] _GEN_770;
  wire [3:0] _GEN_771;
  wire [3:0] _GEN_772;
  wire [3:0] _GEN_773;
  wire [3:0] _GEN_774;
  wire [3:0] _GEN_775;
  wire [3:0] _GEN_776;
  wire [3:0] _GEN_777;
  wire [3:0] _GEN_778;
  wire [3:0] _GEN_779;
  wire [3:0] _GEN_780;
  wire [3:0] _GEN_781;
  wire [3:0] _GEN_782;
  wire [3:0] _GEN_783;
  wire [3:0] _GEN_784;
  wire [3:0] _GEN_785;
  wire [3:0] _GEN_786;
  wire [3:0] _GEN_787;
  wire [3:0] _GEN_788;
  wire [3:0] _GEN_789;
  wire [3:0] _GEN_790;
  wire [3:0] _GEN_791;
  wire [3:0] _GEN_792;
  wire [3:0] _GEN_793;
  wire [3:0] _GEN_794;
  wire [3:0] _GEN_795;
  wire [3:0] _GEN_796;
  wire [3:0] _GEN_797;
  wire [3:0] _GEN_798;
  wire [3:0] _GEN_799;
  wire [3:0] _GEN_800;
  wire [3:0] _GEN_801;
  wire [6:0] _T_212;
  wire [5:0] _T_213;
  wire [3:0] _T_215;
  wire [3:0] _GEN_12;
  wire [3:0] _GEN_802;
  wire [3:0] _GEN_803;
  wire [3:0] _GEN_804;
  wire [3:0] _GEN_805;
  wire [3:0] _GEN_806;
  wire [3:0] _GEN_807;
  wire [3:0] _GEN_808;
  wire [3:0] _GEN_809;
  wire [3:0] _GEN_810;
  wire [3:0] _GEN_811;
  wire [3:0] _GEN_812;
  wire [3:0] _GEN_813;
  wire [3:0] _GEN_814;
  wire [3:0] _GEN_815;
  wire [3:0] _GEN_816;
  wire [3:0] _GEN_817;
  wire [3:0] _GEN_818;
  wire [3:0] _GEN_819;
  wire [3:0] _GEN_820;
  wire [3:0] _GEN_821;
  wire [3:0] _GEN_822;
  wire [3:0] _GEN_823;
  wire [3:0] _GEN_824;
  wire [3:0] _GEN_825;
  wire [3:0] _GEN_826;
  wire [3:0] _GEN_827;
  wire [3:0] _GEN_828;
  wire [3:0] _GEN_829;
  wire [3:0] _GEN_830;
  wire [3:0] _GEN_831;
  wire [3:0] _GEN_832;
  wire [3:0] _GEN_833;
  wire [3:0] _GEN_834;
  wire [3:0] _GEN_835;
  wire [3:0] _GEN_836;
  wire [3:0] _GEN_837;
  wire [3:0] _GEN_838;
  wire [3:0] _GEN_839;
  wire [3:0] _GEN_840;
  wire [3:0] _GEN_841;
  wire [3:0] _GEN_842;
  wire [3:0] _GEN_843;
  wire [3:0] _GEN_844;
  wire [3:0] _GEN_845;
  wire [3:0] _GEN_846;
  wire [3:0] _GEN_847;
  wire [3:0] _GEN_848;
  wire [3:0] _GEN_849;
  wire [3:0] _GEN_850;
  wire [3:0] _GEN_851;
  wire [3:0] _GEN_852;
  wire [3:0] _GEN_853;
  wire [3:0] _GEN_854;
  wire [3:0] _GEN_855;
  wire [3:0] _GEN_856;
  wire [3:0] _GEN_857;
  wire [3:0] _GEN_858;
  wire [3:0] _GEN_859;
  wire [3:0] _GEN_860;
  wire [3:0] _GEN_861;
  wire [3:0] _GEN_862;
  wire [3:0] _GEN_863;
  wire [3:0] _GEN_864;
  wire [3:0] _GEN_865;
  wire [6:0] _T_217;
  wire [5:0] _T_218;
  wire [3:0] _T_220;
  wire [3:0] _GEN_13;
  wire [3:0] _GEN_866;
  wire [3:0] _GEN_867;
  wire [3:0] _GEN_868;
  wire [3:0] _GEN_869;
  wire [3:0] _GEN_870;
  wire [3:0] _GEN_871;
  wire [3:0] _GEN_872;
  wire [3:0] _GEN_873;
  wire [3:0] _GEN_874;
  wire [3:0] _GEN_875;
  wire [3:0] _GEN_876;
  wire [3:0] _GEN_877;
  wire [3:0] _GEN_878;
  wire [3:0] _GEN_879;
  wire [3:0] _GEN_880;
  wire [3:0] _GEN_881;
  wire [3:0] _GEN_882;
  wire [3:0] _GEN_883;
  wire [3:0] _GEN_884;
  wire [3:0] _GEN_885;
  wire [3:0] _GEN_886;
  wire [3:0] _GEN_887;
  wire [3:0] _GEN_888;
  wire [3:0] _GEN_889;
  wire [3:0] _GEN_890;
  wire [3:0] _GEN_891;
  wire [3:0] _GEN_892;
  wire [3:0] _GEN_893;
  wire [3:0] _GEN_894;
  wire [3:0] _GEN_895;
  wire [3:0] _GEN_896;
  wire [3:0] _GEN_897;
  wire [3:0] _GEN_898;
  wire [3:0] _GEN_899;
  wire [3:0] _GEN_900;
  wire [3:0] _GEN_901;
  wire [3:0] _GEN_902;
  wire [3:0] _GEN_903;
  wire [3:0] _GEN_904;
  wire [3:0] _GEN_905;
  wire [3:0] _GEN_906;
  wire [3:0] _GEN_907;
  wire [3:0] _GEN_908;
  wire [3:0] _GEN_909;
  wire [3:0] _GEN_910;
  wire [3:0] _GEN_911;
  wire [3:0] _GEN_912;
  wire [3:0] _GEN_913;
  wire [3:0] _GEN_914;
  wire [3:0] _GEN_915;
  wire [3:0] _GEN_916;
  wire [3:0] _GEN_917;
  wire [3:0] _GEN_918;
  wire [3:0] _GEN_919;
  wire [3:0] _GEN_920;
  wire [3:0] _GEN_921;
  wire [3:0] _GEN_922;
  wire [3:0] _GEN_923;
  wire [3:0] _GEN_924;
  wire [3:0] _GEN_925;
  wire [3:0] _GEN_926;
  wire [3:0] _GEN_927;
  wire [3:0] _GEN_928;
  wire [3:0] _GEN_929;
  wire [6:0] _T_222;
  wire [5:0] _T_223;
  wire [3:0] _T_225;
  wire [3:0] _GEN_14;
  wire [3:0] _GEN_930;
  wire [3:0] _GEN_931;
  wire [3:0] _GEN_932;
  wire [3:0] _GEN_933;
  wire [3:0] _GEN_934;
  wire [3:0] _GEN_935;
  wire [3:0] _GEN_936;
  wire [3:0] _GEN_937;
  wire [3:0] _GEN_938;
  wire [3:0] _GEN_939;
  wire [3:0] _GEN_940;
  wire [3:0] _GEN_941;
  wire [3:0] _GEN_942;
  wire [3:0] _GEN_943;
  wire [3:0] _GEN_944;
  wire [3:0] _GEN_945;
  wire [3:0] _GEN_946;
  wire [3:0] _GEN_947;
  wire [3:0] _GEN_948;
  wire [3:0] _GEN_949;
  wire [3:0] _GEN_950;
  wire [3:0] _GEN_951;
  wire [3:0] _GEN_952;
  wire [3:0] _GEN_953;
  wire [3:0] _GEN_954;
  wire [3:0] _GEN_955;
  wire [3:0] _GEN_956;
  wire [3:0] _GEN_957;
  wire [3:0] _GEN_958;
  wire [3:0] _GEN_959;
  wire [3:0] _GEN_960;
  wire [3:0] _GEN_961;
  wire [3:0] _GEN_962;
  wire [3:0] _GEN_963;
  wire [3:0] _GEN_964;
  wire [3:0] _GEN_965;
  wire [3:0] _GEN_966;
  wire [3:0] _GEN_967;
  wire [3:0] _GEN_968;
  wire [3:0] _GEN_969;
  wire [3:0] _GEN_970;
  wire [3:0] _GEN_971;
  wire [3:0] _GEN_972;
  wire [3:0] _GEN_973;
  wire [3:0] _GEN_974;
  wire [3:0] _GEN_975;
  wire [3:0] _GEN_976;
  wire [3:0] _GEN_977;
  wire [3:0] _GEN_978;
  wire [3:0] _GEN_979;
  wire [3:0] _GEN_980;
  wire [3:0] _GEN_981;
  wire [3:0] _GEN_982;
  wire [3:0] _GEN_983;
  wire [3:0] _GEN_984;
  wire [3:0] _GEN_985;
  wire [3:0] _GEN_986;
  wire [3:0] _GEN_987;
  wire [3:0] _GEN_988;
  wire [3:0] _GEN_989;
  wire [3:0] _GEN_990;
  wire [3:0] _GEN_991;
  wire [3:0] _GEN_992;
  wire [3:0] _GEN_993;
  wire [6:0] _T_227;
  wire [5:0] _T_228;
  wire [3:0] _T_230;
  wire [3:0] _GEN_15;
  wire [3:0] _GEN_994;
  wire [3:0] _GEN_995;
  wire [3:0] _GEN_996;
  wire [3:0] _GEN_997;
  wire [3:0] _GEN_998;
  wire [3:0] _GEN_999;
  wire [3:0] _GEN_1000;
  wire [3:0] _GEN_1001;
  wire [3:0] _GEN_1002;
  wire [3:0] _GEN_1003;
  wire [3:0] _GEN_1004;
  wire [3:0] _GEN_1005;
  wire [3:0] _GEN_1006;
  wire [3:0] _GEN_1007;
  wire [3:0] _GEN_1008;
  wire [3:0] _GEN_1009;
  wire [3:0] _GEN_1010;
  wire [3:0] _GEN_1011;
  wire [3:0] _GEN_1012;
  wire [3:0] _GEN_1013;
  wire [3:0] _GEN_1014;
  wire [3:0] _GEN_1015;
  wire [3:0] _GEN_1016;
  wire [3:0] _GEN_1017;
  wire [3:0] _GEN_1018;
  wire [3:0] _GEN_1019;
  wire [3:0] _GEN_1020;
  wire [3:0] _GEN_1021;
  wire [3:0] _GEN_1022;
  wire [3:0] _GEN_1023;
  wire [3:0] _GEN_1024;
  wire [3:0] _GEN_1025;
  wire [3:0] _GEN_1026;
  wire [3:0] _GEN_1027;
  wire [3:0] _GEN_1028;
  wire [3:0] _GEN_1029;
  wire [3:0] _GEN_1030;
  wire [3:0] _GEN_1031;
  wire [3:0] _GEN_1032;
  wire [3:0] _GEN_1033;
  wire [3:0] _GEN_1034;
  wire [3:0] _GEN_1035;
  wire [3:0] _GEN_1036;
  wire [3:0] _GEN_1037;
  wire [3:0] _GEN_1038;
  wire [3:0] _GEN_1039;
  wire [3:0] _GEN_1040;
  wire [3:0] _GEN_1041;
  wire [3:0] _GEN_1042;
  wire [3:0] _GEN_1043;
  wire [3:0] _GEN_1044;
  wire [3:0] _GEN_1045;
  wire [3:0] _GEN_1046;
  wire [3:0] _GEN_1047;
  wire [3:0] _GEN_1048;
  wire [3:0] _GEN_1049;
  wire [3:0] _GEN_1050;
  wire [3:0] _GEN_1051;
  wire [3:0] _GEN_1052;
  wire [3:0] _GEN_1053;
  wire [3:0] _GEN_1054;
  wire [3:0] _GEN_1055;
  wire [3:0] _GEN_1056;
  wire [3:0] _GEN_1057;
  wire [6:0] _T_232;
  wire [5:0] _T_233;
  wire [3:0] _T_235;
  wire [3:0] _GEN_16;
  wire [3:0] _GEN_1058;
  wire [3:0] _GEN_1059;
  wire [3:0] _GEN_1060;
  wire [3:0] _GEN_1061;
  wire [3:0] _GEN_1062;
  wire [3:0] _GEN_1063;
  wire [3:0] _GEN_1064;
  wire [3:0] _GEN_1065;
  wire [3:0] _GEN_1066;
  wire [3:0] _GEN_1067;
  wire [3:0] _GEN_1068;
  wire [3:0] _GEN_1069;
  wire [3:0] _GEN_1070;
  wire [3:0] _GEN_1071;
  wire [3:0] _GEN_1072;
  wire [3:0] _GEN_1073;
  wire [3:0] _GEN_1074;
  wire [3:0] _GEN_1075;
  wire [3:0] _GEN_1076;
  wire [3:0] _GEN_1077;
  wire [3:0] _GEN_1078;
  wire [3:0] _GEN_1079;
  wire [3:0] _GEN_1080;
  wire [3:0] _GEN_1081;
  wire [3:0] _GEN_1082;
  wire [3:0] _GEN_1083;
  wire [3:0] _GEN_1084;
  wire [3:0] _GEN_1085;
  wire [3:0] _GEN_1086;
  wire [3:0] _GEN_1087;
  wire [3:0] _GEN_1088;
  wire [3:0] _GEN_1089;
  wire [3:0] _GEN_1090;
  wire [3:0] _GEN_1091;
  wire [3:0] _GEN_1092;
  wire [3:0] _GEN_1093;
  wire [3:0] _GEN_1094;
  wire [3:0] _GEN_1095;
  wire [3:0] _GEN_1096;
  wire [3:0] _GEN_1097;
  wire [3:0] _GEN_1098;
  wire [3:0] _GEN_1099;
  wire [3:0] _GEN_1100;
  wire [3:0] _GEN_1101;
  wire [3:0] _GEN_1102;
  wire [3:0] _GEN_1103;
  wire [3:0] _GEN_1104;
  wire [3:0] _GEN_1105;
  wire [3:0] _GEN_1106;
  wire [3:0] _GEN_1107;
  wire [3:0] _GEN_1108;
  wire [3:0] _GEN_1109;
  wire [3:0] _GEN_1110;
  wire [3:0] _GEN_1111;
  wire [3:0] _GEN_1112;
  wire [3:0] _GEN_1113;
  wire [3:0] _GEN_1114;
  wire [3:0] _GEN_1115;
  wire [3:0] _GEN_1116;
  wire [3:0] _GEN_1117;
  wire [3:0] _GEN_1118;
  wire [3:0] _GEN_1119;
  wire [3:0] _GEN_1120;
  wire [3:0] _GEN_1121;
  wire [6:0] _T_237;
  wire [5:0] _T_238;
  wire [3:0] _T_240;
  wire [3:0] _GEN_17;
  wire [3:0] _GEN_1122;
  wire [3:0] _GEN_1123;
  wire [3:0] _GEN_1124;
  wire [3:0] _GEN_1125;
  wire [3:0] _GEN_1126;
  wire [3:0] _GEN_1127;
  wire [3:0] _GEN_1128;
  wire [3:0] _GEN_1129;
  wire [3:0] _GEN_1130;
  wire [3:0] _GEN_1131;
  wire [3:0] _GEN_1132;
  wire [3:0] _GEN_1133;
  wire [3:0] _GEN_1134;
  wire [3:0] _GEN_1135;
  wire [3:0] _GEN_1136;
  wire [3:0] _GEN_1137;
  wire [3:0] _GEN_1138;
  wire [3:0] _GEN_1139;
  wire [3:0] _GEN_1140;
  wire [3:0] _GEN_1141;
  wire [3:0] _GEN_1142;
  wire [3:0] _GEN_1143;
  wire [3:0] _GEN_1144;
  wire [3:0] _GEN_1145;
  wire [3:0] _GEN_1146;
  wire [3:0] _GEN_1147;
  wire [3:0] _GEN_1148;
  wire [3:0] _GEN_1149;
  wire [3:0] _GEN_1150;
  wire [3:0] _GEN_1151;
  wire [3:0] _GEN_1152;
  wire [3:0] _GEN_1153;
  wire [3:0] _GEN_1154;
  wire [3:0] _GEN_1155;
  wire [3:0] _GEN_1156;
  wire [3:0] _GEN_1157;
  wire [3:0] _GEN_1158;
  wire [3:0] _GEN_1159;
  wire [3:0] _GEN_1160;
  wire [3:0] _GEN_1161;
  wire [3:0] _GEN_1162;
  wire [3:0] _GEN_1163;
  wire [3:0] _GEN_1164;
  wire [3:0] _GEN_1165;
  wire [3:0] _GEN_1166;
  wire [3:0] _GEN_1167;
  wire [3:0] _GEN_1168;
  wire [3:0] _GEN_1169;
  wire [3:0] _GEN_1170;
  wire [3:0] _GEN_1171;
  wire [3:0] _GEN_1172;
  wire [3:0] _GEN_1173;
  wire [3:0] _GEN_1174;
  wire [3:0] _GEN_1175;
  wire [3:0] _GEN_1176;
  wire [3:0] _GEN_1177;
  wire [3:0] _GEN_1178;
  wire [3:0] _GEN_1179;
  wire [3:0] _GEN_1180;
  wire [3:0] _GEN_1181;
  wire [3:0] _GEN_1182;
  wire [3:0] _GEN_1183;
  wire [3:0] _GEN_1184;
  wire [3:0] _GEN_1185;
  wire [6:0] _T_242;
  wire [5:0] _T_243;
  wire [3:0] _T_245;
  wire [3:0] _GEN_18;
  wire [3:0] _GEN_1186;
  wire [3:0] _GEN_1187;
  wire [3:0] _GEN_1188;
  wire [3:0] _GEN_1189;
  wire [3:0] _GEN_1190;
  wire [3:0] _GEN_1191;
  wire [3:0] _GEN_1192;
  wire [3:0] _GEN_1193;
  wire [3:0] _GEN_1194;
  wire [3:0] _GEN_1195;
  wire [3:0] _GEN_1196;
  wire [3:0] _GEN_1197;
  wire [3:0] _GEN_1198;
  wire [3:0] _GEN_1199;
  wire [3:0] _GEN_1200;
  wire [3:0] _GEN_1201;
  wire [3:0] _GEN_1202;
  wire [3:0] _GEN_1203;
  wire [3:0] _GEN_1204;
  wire [3:0] _GEN_1205;
  wire [3:0] _GEN_1206;
  wire [3:0] _GEN_1207;
  wire [3:0] _GEN_1208;
  wire [3:0] _GEN_1209;
  wire [3:0] _GEN_1210;
  wire [3:0] _GEN_1211;
  wire [3:0] _GEN_1212;
  wire [3:0] _GEN_1213;
  wire [3:0] _GEN_1214;
  wire [3:0] _GEN_1215;
  wire [3:0] _GEN_1216;
  wire [3:0] _GEN_1217;
  wire [3:0] _GEN_1218;
  wire [3:0] _GEN_1219;
  wire [3:0] _GEN_1220;
  wire [3:0] _GEN_1221;
  wire [3:0] _GEN_1222;
  wire [3:0] _GEN_1223;
  wire [3:0] _GEN_1224;
  wire [3:0] _GEN_1225;
  wire [3:0] _GEN_1226;
  wire [3:0] _GEN_1227;
  wire [3:0] _GEN_1228;
  wire [3:0] _GEN_1229;
  wire [3:0] _GEN_1230;
  wire [3:0] _GEN_1231;
  wire [3:0] _GEN_1232;
  wire [3:0] _GEN_1233;
  wire [3:0] _GEN_1234;
  wire [3:0] _GEN_1235;
  wire [3:0] _GEN_1236;
  wire [3:0] _GEN_1237;
  wire [3:0] _GEN_1238;
  wire [3:0] _GEN_1239;
  wire [3:0] _GEN_1240;
  wire [3:0] _GEN_1241;
  wire [3:0] _GEN_1242;
  wire [3:0] _GEN_1243;
  wire [3:0] _GEN_1244;
  wire [3:0] _GEN_1245;
  wire [3:0] _GEN_1246;
  wire [3:0] _GEN_1247;
  wire [3:0] _GEN_1248;
  wire [3:0] _GEN_1249;
  wire [6:0] _T_247;
  wire [5:0] _T_248;
  wire [3:0] _T_250;
  wire [3:0] _GEN_19;
  wire [3:0] _GEN_1250;
  wire [3:0] _GEN_1251;
  wire [3:0] _GEN_1252;
  wire [3:0] _GEN_1253;
  wire [3:0] _GEN_1254;
  wire [3:0] _GEN_1255;
  wire [3:0] _GEN_1256;
  wire [3:0] _GEN_1257;
  wire [3:0] _GEN_1258;
  wire [3:0] _GEN_1259;
  wire [3:0] _GEN_1260;
  wire [3:0] _GEN_1261;
  wire [3:0] _GEN_1262;
  wire [3:0] _GEN_1263;
  wire [3:0] _GEN_1264;
  wire [3:0] _GEN_1265;
  wire [3:0] _GEN_1266;
  wire [3:0] _GEN_1267;
  wire [3:0] _GEN_1268;
  wire [3:0] _GEN_1269;
  wire [3:0] _GEN_1270;
  wire [3:0] _GEN_1271;
  wire [3:0] _GEN_1272;
  wire [3:0] _GEN_1273;
  wire [3:0] _GEN_1274;
  wire [3:0] _GEN_1275;
  wire [3:0] _GEN_1276;
  wire [3:0] _GEN_1277;
  wire [3:0] _GEN_1278;
  wire [3:0] _GEN_1279;
  wire [3:0] _GEN_1280;
  wire [3:0] _GEN_1281;
  wire [3:0] _GEN_1282;
  wire [3:0] _GEN_1283;
  wire [3:0] _GEN_1284;
  wire [3:0] _GEN_1285;
  wire [3:0] _GEN_1286;
  wire [3:0] _GEN_1287;
  wire [3:0] _GEN_1288;
  wire [3:0] _GEN_1289;
  wire [3:0] _GEN_1290;
  wire [3:0] _GEN_1291;
  wire [3:0] _GEN_1292;
  wire [3:0] _GEN_1293;
  wire [3:0] _GEN_1294;
  wire [3:0] _GEN_1295;
  wire [3:0] _GEN_1296;
  wire [3:0] _GEN_1297;
  wire [3:0] _GEN_1298;
  wire [3:0] _GEN_1299;
  wire [3:0] _GEN_1300;
  wire [3:0] _GEN_1301;
  wire [3:0] _GEN_1302;
  wire [3:0] _GEN_1303;
  wire [3:0] _GEN_1304;
  wire [3:0] _GEN_1305;
  wire [3:0] _GEN_1306;
  wire [3:0] _GEN_1307;
  wire [3:0] _GEN_1308;
  wire [3:0] _GEN_1309;
  wire [3:0] _GEN_1310;
  wire [3:0] _GEN_1311;
  wire [3:0] _GEN_1312;
  wire [3:0] _GEN_1313;
  wire [6:0] _T_252;
  wire [5:0] _T_253;
  wire [3:0] _T_255;
  wire [3:0] _GEN_20;
  wire [3:0] _GEN_1314;
  wire [3:0] _GEN_1315;
  wire [3:0] _GEN_1316;
  wire [3:0] _GEN_1317;
  wire [3:0] _GEN_1318;
  wire [3:0] _GEN_1319;
  wire [3:0] _GEN_1320;
  wire [3:0] _GEN_1321;
  wire [3:0] _GEN_1322;
  wire [3:0] _GEN_1323;
  wire [3:0] _GEN_1324;
  wire [3:0] _GEN_1325;
  wire [3:0] _GEN_1326;
  wire [3:0] _GEN_1327;
  wire [3:0] _GEN_1328;
  wire [3:0] _GEN_1329;
  wire [3:0] _GEN_1330;
  wire [3:0] _GEN_1331;
  wire [3:0] _GEN_1332;
  wire [3:0] _GEN_1333;
  wire [3:0] _GEN_1334;
  wire [3:0] _GEN_1335;
  wire [3:0] _GEN_1336;
  wire [3:0] _GEN_1337;
  wire [3:0] _GEN_1338;
  wire [3:0] _GEN_1339;
  wire [3:0] _GEN_1340;
  wire [3:0] _GEN_1341;
  wire [3:0] _GEN_1342;
  wire [3:0] _GEN_1343;
  wire [3:0] _GEN_1344;
  wire [3:0] _GEN_1345;
  wire [3:0] _GEN_1346;
  wire [3:0] _GEN_1347;
  wire [3:0] _GEN_1348;
  wire [3:0] _GEN_1349;
  wire [3:0] _GEN_1350;
  wire [3:0] _GEN_1351;
  wire [3:0] _GEN_1352;
  wire [3:0] _GEN_1353;
  wire [3:0] _GEN_1354;
  wire [3:0] _GEN_1355;
  wire [3:0] _GEN_1356;
  wire [3:0] _GEN_1357;
  wire [3:0] _GEN_1358;
  wire [3:0] _GEN_1359;
  wire [3:0] _GEN_1360;
  wire [3:0] _GEN_1361;
  wire [3:0] _GEN_1362;
  wire [3:0] _GEN_1363;
  wire [3:0] _GEN_1364;
  wire [3:0] _GEN_1365;
  wire [3:0] _GEN_1366;
  wire [3:0] _GEN_1367;
  wire [3:0] _GEN_1368;
  wire [3:0] _GEN_1369;
  wire [3:0] _GEN_1370;
  wire [3:0] _GEN_1371;
  wire [3:0] _GEN_1372;
  wire [3:0] _GEN_1373;
  wire [3:0] _GEN_1374;
  wire [3:0] _GEN_1375;
  wire [3:0] _GEN_1376;
  wire [3:0] _GEN_1377;
  wire [6:0] _T_257;
  wire [5:0] _T_258;
  wire [3:0] _T_260;
  wire [3:0] _GEN_21;
  wire [3:0] _GEN_1378;
  wire [3:0] _GEN_1379;
  wire [3:0] _GEN_1380;
  wire [3:0] _GEN_1381;
  wire [3:0] _GEN_1382;
  wire [3:0] _GEN_1383;
  wire [3:0] _GEN_1384;
  wire [3:0] _GEN_1385;
  wire [3:0] _GEN_1386;
  wire [3:0] _GEN_1387;
  wire [3:0] _GEN_1388;
  wire [3:0] _GEN_1389;
  wire [3:0] _GEN_1390;
  wire [3:0] _GEN_1391;
  wire [3:0] _GEN_1392;
  wire [3:0] _GEN_1393;
  wire [3:0] _GEN_1394;
  wire [3:0] _GEN_1395;
  wire [3:0] _GEN_1396;
  wire [3:0] _GEN_1397;
  wire [3:0] _GEN_1398;
  wire [3:0] _GEN_1399;
  wire [3:0] _GEN_1400;
  wire [3:0] _GEN_1401;
  wire [3:0] _GEN_1402;
  wire [3:0] _GEN_1403;
  wire [3:0] _GEN_1404;
  wire [3:0] _GEN_1405;
  wire [3:0] _GEN_1406;
  wire [3:0] _GEN_1407;
  wire [3:0] _GEN_1408;
  wire [3:0] _GEN_1409;
  wire [3:0] _GEN_1410;
  wire [3:0] _GEN_1411;
  wire [3:0] _GEN_1412;
  wire [3:0] _GEN_1413;
  wire [3:0] _GEN_1414;
  wire [3:0] _GEN_1415;
  wire [3:0] _GEN_1416;
  wire [3:0] _GEN_1417;
  wire [3:0] _GEN_1418;
  wire [3:0] _GEN_1419;
  wire [3:0] _GEN_1420;
  wire [3:0] _GEN_1421;
  wire [3:0] _GEN_1422;
  wire [3:0] _GEN_1423;
  wire [3:0] _GEN_1424;
  wire [3:0] _GEN_1425;
  wire [3:0] _GEN_1426;
  wire [3:0] _GEN_1427;
  wire [3:0] _GEN_1428;
  wire [3:0] _GEN_1429;
  wire [3:0] _GEN_1430;
  wire [3:0] _GEN_1431;
  wire [3:0] _GEN_1432;
  wire [3:0] _GEN_1433;
  wire [3:0] _GEN_1434;
  wire [3:0] _GEN_1435;
  wire [3:0] _GEN_1436;
  wire [3:0] _GEN_1437;
  wire [3:0] _GEN_1438;
  wire [3:0] _GEN_1439;
  wire [3:0] _GEN_1440;
  wire [3:0] _GEN_1441;
  wire [6:0] _T_262;
  wire [5:0] _T_263;
  wire [3:0] _T_265;
  wire [3:0] _GEN_22;
  wire [3:0] _GEN_1442;
  wire [3:0] _GEN_1443;
  wire [3:0] _GEN_1444;
  wire [3:0] _GEN_1445;
  wire [3:0] _GEN_1446;
  wire [3:0] _GEN_1447;
  wire [3:0] _GEN_1448;
  wire [3:0] _GEN_1449;
  wire [3:0] _GEN_1450;
  wire [3:0] _GEN_1451;
  wire [3:0] _GEN_1452;
  wire [3:0] _GEN_1453;
  wire [3:0] _GEN_1454;
  wire [3:0] _GEN_1455;
  wire [3:0] _GEN_1456;
  wire [3:0] _GEN_1457;
  wire [3:0] _GEN_1458;
  wire [3:0] _GEN_1459;
  wire [3:0] _GEN_1460;
  wire [3:0] _GEN_1461;
  wire [3:0] _GEN_1462;
  wire [3:0] _GEN_1463;
  wire [3:0] _GEN_1464;
  wire [3:0] _GEN_1465;
  wire [3:0] _GEN_1466;
  wire [3:0] _GEN_1467;
  wire [3:0] _GEN_1468;
  wire [3:0] _GEN_1469;
  wire [3:0] _GEN_1470;
  wire [3:0] _GEN_1471;
  wire [3:0] _GEN_1472;
  wire [3:0] _GEN_1473;
  wire [3:0] _GEN_1474;
  wire [3:0] _GEN_1475;
  wire [3:0] _GEN_1476;
  wire [3:0] _GEN_1477;
  wire [3:0] _GEN_1478;
  wire [3:0] _GEN_1479;
  wire [3:0] _GEN_1480;
  wire [3:0] _GEN_1481;
  wire [3:0] _GEN_1482;
  wire [3:0] _GEN_1483;
  wire [3:0] _GEN_1484;
  wire [3:0] _GEN_1485;
  wire [3:0] _GEN_1486;
  wire [3:0] _GEN_1487;
  wire [3:0] _GEN_1488;
  wire [3:0] _GEN_1489;
  wire [3:0] _GEN_1490;
  wire [3:0] _GEN_1491;
  wire [3:0] _GEN_1492;
  wire [3:0] _GEN_1493;
  wire [3:0] _GEN_1494;
  wire [3:0] _GEN_1495;
  wire [3:0] _GEN_1496;
  wire [3:0] _GEN_1497;
  wire [3:0] _GEN_1498;
  wire [3:0] _GEN_1499;
  wire [3:0] _GEN_1500;
  wire [3:0] _GEN_1501;
  wire [3:0] _GEN_1502;
  wire [3:0] _GEN_1503;
  wire [3:0] _GEN_1504;
  wire [3:0] _GEN_1505;
  wire [6:0] _T_267;
  wire [5:0] _T_268;
  wire [3:0] _T_270;
  wire [3:0] _GEN_23;
  wire [3:0] _GEN_1506;
  wire [3:0] _GEN_1507;
  wire [3:0] _GEN_1508;
  wire [3:0] _GEN_1509;
  wire [3:0] _GEN_1510;
  wire [3:0] _GEN_1511;
  wire [3:0] _GEN_1512;
  wire [3:0] _GEN_1513;
  wire [3:0] _GEN_1514;
  wire [3:0] _GEN_1515;
  wire [3:0] _GEN_1516;
  wire [3:0] _GEN_1517;
  wire [3:0] _GEN_1518;
  wire [3:0] _GEN_1519;
  wire [3:0] _GEN_1520;
  wire [3:0] _GEN_1521;
  wire [3:0] _GEN_1522;
  wire [3:0] _GEN_1523;
  wire [3:0] _GEN_1524;
  wire [3:0] _GEN_1525;
  wire [3:0] _GEN_1526;
  wire [3:0] _GEN_1527;
  wire [3:0] _GEN_1528;
  wire [3:0] _GEN_1529;
  wire [3:0] _GEN_1530;
  wire [3:0] _GEN_1531;
  wire [3:0] _GEN_1532;
  wire [3:0] _GEN_1533;
  wire [3:0] _GEN_1534;
  wire [3:0] _GEN_1535;
  wire [3:0] _GEN_1536;
  wire [3:0] _GEN_1537;
  wire [3:0] _GEN_1538;
  wire [3:0] _GEN_1539;
  wire [3:0] _GEN_1540;
  wire [3:0] _GEN_1541;
  wire [3:0] _GEN_1542;
  wire [3:0] _GEN_1543;
  wire [3:0] _GEN_1544;
  wire [3:0] _GEN_1545;
  wire [3:0] _GEN_1546;
  wire [3:0] _GEN_1547;
  wire [3:0] _GEN_1548;
  wire [3:0] _GEN_1549;
  wire [3:0] _GEN_1550;
  wire [3:0] _GEN_1551;
  wire [3:0] _GEN_1552;
  wire [3:0] _GEN_1553;
  wire [3:0] _GEN_1554;
  wire [3:0] _GEN_1555;
  wire [3:0] _GEN_1556;
  wire [3:0] _GEN_1557;
  wire [3:0] _GEN_1558;
  wire [3:0] _GEN_1559;
  wire [3:0] _GEN_1560;
  wire [3:0] _GEN_1561;
  wire [3:0] _GEN_1562;
  wire [3:0] _GEN_1563;
  wire [3:0] _GEN_1564;
  wire [3:0] _GEN_1565;
  wire [3:0] _GEN_1566;
  wire [3:0] _GEN_1567;
  wire [3:0] _GEN_1568;
  wire [3:0] _GEN_1569;
  wire [6:0] _T_272;
  wire [5:0] _T_273;
  wire [3:0] _T_275;
  wire [3:0] _GEN_24;
  wire [3:0] _GEN_1570;
  wire [3:0] _GEN_1571;
  wire [3:0] _GEN_1572;
  wire [3:0] _GEN_1573;
  wire [3:0] _GEN_1574;
  wire [3:0] _GEN_1575;
  wire [3:0] _GEN_1576;
  wire [3:0] _GEN_1577;
  wire [3:0] _GEN_1578;
  wire [3:0] _GEN_1579;
  wire [3:0] _GEN_1580;
  wire [3:0] _GEN_1581;
  wire [3:0] _GEN_1582;
  wire [3:0] _GEN_1583;
  wire [3:0] _GEN_1584;
  wire [3:0] _GEN_1585;
  wire [3:0] _GEN_1586;
  wire [3:0] _GEN_1587;
  wire [3:0] _GEN_1588;
  wire [3:0] _GEN_1589;
  wire [3:0] _GEN_1590;
  wire [3:0] _GEN_1591;
  wire [3:0] _GEN_1592;
  wire [3:0] _GEN_1593;
  wire [3:0] _GEN_1594;
  wire [3:0] _GEN_1595;
  wire [3:0] _GEN_1596;
  wire [3:0] _GEN_1597;
  wire [3:0] _GEN_1598;
  wire [3:0] _GEN_1599;
  wire [3:0] _GEN_1600;
  wire [3:0] _GEN_1601;
  wire [3:0] _GEN_1602;
  wire [3:0] _GEN_1603;
  wire [3:0] _GEN_1604;
  wire [3:0] _GEN_1605;
  wire [3:0] _GEN_1606;
  wire [3:0] _GEN_1607;
  wire [3:0] _GEN_1608;
  wire [3:0] _GEN_1609;
  wire [3:0] _GEN_1610;
  wire [3:0] _GEN_1611;
  wire [3:0] _GEN_1612;
  wire [3:0] _GEN_1613;
  wire [3:0] _GEN_1614;
  wire [3:0] _GEN_1615;
  wire [3:0] _GEN_1616;
  wire [3:0] _GEN_1617;
  wire [3:0] _GEN_1618;
  wire [3:0] _GEN_1619;
  wire [3:0] _GEN_1620;
  wire [3:0] _GEN_1621;
  wire [3:0] _GEN_1622;
  wire [3:0] _GEN_1623;
  wire [3:0] _GEN_1624;
  wire [3:0] _GEN_1625;
  wire [3:0] _GEN_1626;
  wire [3:0] _GEN_1627;
  wire [3:0] _GEN_1628;
  wire [3:0] _GEN_1629;
  wire [3:0] _GEN_1630;
  wire [3:0] _GEN_1631;
  wire [3:0] _GEN_1632;
  wire [3:0] _GEN_1633;
  wire [6:0] _T_277;
  wire [5:0] _T_278;
  wire [3:0] _T_280;
  wire [3:0] _GEN_25;
  wire [3:0] _GEN_1634;
  wire [3:0] _GEN_1635;
  wire [3:0] _GEN_1636;
  wire [3:0] _GEN_1637;
  wire [3:0] _GEN_1638;
  wire [3:0] _GEN_1639;
  wire [3:0] _GEN_1640;
  wire [3:0] _GEN_1641;
  wire [3:0] _GEN_1642;
  wire [3:0] _GEN_1643;
  wire [3:0] _GEN_1644;
  wire [3:0] _GEN_1645;
  wire [3:0] _GEN_1646;
  wire [3:0] _GEN_1647;
  wire [3:0] _GEN_1648;
  wire [3:0] _GEN_1649;
  wire [3:0] _GEN_1650;
  wire [3:0] _GEN_1651;
  wire [3:0] _GEN_1652;
  wire [3:0] _GEN_1653;
  wire [3:0] _GEN_1654;
  wire [3:0] _GEN_1655;
  wire [3:0] _GEN_1656;
  wire [3:0] _GEN_1657;
  wire [3:0] _GEN_1658;
  wire [3:0] _GEN_1659;
  wire [3:0] _GEN_1660;
  wire [3:0] _GEN_1661;
  wire [3:0] _GEN_1662;
  wire [3:0] _GEN_1663;
  wire [3:0] _GEN_1664;
  wire [3:0] _GEN_1665;
  wire [3:0] _GEN_1666;
  wire [3:0] _GEN_1667;
  wire [3:0] _GEN_1668;
  wire [3:0] _GEN_1669;
  wire [3:0] _GEN_1670;
  wire [3:0] _GEN_1671;
  wire [3:0] _GEN_1672;
  wire [3:0] _GEN_1673;
  wire [3:0] _GEN_1674;
  wire [3:0] _GEN_1675;
  wire [3:0] _GEN_1676;
  wire [3:0] _GEN_1677;
  wire [3:0] _GEN_1678;
  wire [3:0] _GEN_1679;
  wire [3:0] _GEN_1680;
  wire [3:0] _GEN_1681;
  wire [3:0] _GEN_1682;
  wire [3:0] _GEN_1683;
  wire [3:0] _GEN_1684;
  wire [3:0] _GEN_1685;
  wire [3:0] _GEN_1686;
  wire [3:0] _GEN_1687;
  wire [3:0] _GEN_1688;
  wire [3:0] _GEN_1689;
  wire [3:0] _GEN_1690;
  wire [3:0] _GEN_1691;
  wire [3:0] _GEN_1692;
  wire [3:0] _GEN_1693;
  wire [3:0] _GEN_1694;
  wire [3:0] _GEN_1695;
  wire [3:0] _GEN_1696;
  wire [3:0] _GEN_1697;
  wire [6:0] _T_282;
  wire [5:0] _T_283;
  wire [3:0] _T_285;
  wire [3:0] _GEN_26;
  wire [3:0] _GEN_1698;
  wire [3:0] _GEN_1699;
  wire [3:0] _GEN_1700;
  wire [3:0] _GEN_1701;
  wire [3:0] _GEN_1702;
  wire [3:0] _GEN_1703;
  wire [3:0] _GEN_1704;
  wire [3:0] _GEN_1705;
  wire [3:0] _GEN_1706;
  wire [3:0] _GEN_1707;
  wire [3:0] _GEN_1708;
  wire [3:0] _GEN_1709;
  wire [3:0] _GEN_1710;
  wire [3:0] _GEN_1711;
  wire [3:0] _GEN_1712;
  wire [3:0] _GEN_1713;
  wire [3:0] _GEN_1714;
  wire [3:0] _GEN_1715;
  wire [3:0] _GEN_1716;
  wire [3:0] _GEN_1717;
  wire [3:0] _GEN_1718;
  wire [3:0] _GEN_1719;
  wire [3:0] _GEN_1720;
  wire [3:0] _GEN_1721;
  wire [3:0] _GEN_1722;
  wire [3:0] _GEN_1723;
  wire [3:0] _GEN_1724;
  wire [3:0] _GEN_1725;
  wire [3:0] _GEN_1726;
  wire [3:0] _GEN_1727;
  wire [3:0] _GEN_1728;
  wire [3:0] _GEN_1729;
  wire [3:0] _GEN_1730;
  wire [3:0] _GEN_1731;
  wire [3:0] _GEN_1732;
  wire [3:0] _GEN_1733;
  wire [3:0] _GEN_1734;
  wire [3:0] _GEN_1735;
  wire [3:0] _GEN_1736;
  wire [3:0] _GEN_1737;
  wire [3:0] _GEN_1738;
  wire [3:0] _GEN_1739;
  wire [3:0] _GEN_1740;
  wire [3:0] _GEN_1741;
  wire [3:0] _GEN_1742;
  wire [3:0] _GEN_1743;
  wire [3:0] _GEN_1744;
  wire [3:0] _GEN_1745;
  wire [3:0] _GEN_1746;
  wire [3:0] _GEN_1747;
  wire [3:0] _GEN_1748;
  wire [3:0] _GEN_1749;
  wire [3:0] _GEN_1750;
  wire [3:0] _GEN_1751;
  wire [3:0] _GEN_1752;
  wire [3:0] _GEN_1753;
  wire [3:0] _GEN_1754;
  wire [3:0] _GEN_1755;
  wire [3:0] _GEN_1756;
  wire [3:0] _GEN_1757;
  wire [3:0] _GEN_1758;
  wire [3:0] _GEN_1759;
  wire [3:0] _GEN_1760;
  wire [3:0] _GEN_1761;
  wire [6:0] _T_287;
  wire [5:0] _T_288;
  wire [3:0] _T_290;
  wire [3:0] _GEN_27;
  wire [3:0] _GEN_1762;
  wire [3:0] _GEN_1763;
  wire [3:0] _GEN_1764;
  wire [3:0] _GEN_1765;
  wire [3:0] _GEN_1766;
  wire [3:0] _GEN_1767;
  wire [3:0] _GEN_1768;
  wire [3:0] _GEN_1769;
  wire [3:0] _GEN_1770;
  wire [3:0] _GEN_1771;
  wire [3:0] _GEN_1772;
  wire [3:0] _GEN_1773;
  wire [3:0] _GEN_1774;
  wire [3:0] _GEN_1775;
  wire [3:0] _GEN_1776;
  wire [3:0] _GEN_1777;
  wire [3:0] _GEN_1778;
  wire [3:0] _GEN_1779;
  wire [3:0] _GEN_1780;
  wire [3:0] _GEN_1781;
  wire [3:0] _GEN_1782;
  wire [3:0] _GEN_1783;
  wire [3:0] _GEN_1784;
  wire [3:0] _GEN_1785;
  wire [3:0] _GEN_1786;
  wire [3:0] _GEN_1787;
  wire [3:0] _GEN_1788;
  wire [3:0] _GEN_1789;
  wire [3:0] _GEN_1790;
  wire [3:0] _GEN_1791;
  wire [3:0] _GEN_1792;
  wire [3:0] _GEN_1793;
  wire [3:0] _GEN_1794;
  wire [3:0] _GEN_1795;
  wire [3:0] _GEN_1796;
  wire [3:0] _GEN_1797;
  wire [3:0] _GEN_1798;
  wire [3:0] _GEN_1799;
  wire [3:0] _GEN_1800;
  wire [3:0] _GEN_1801;
  wire [3:0] _GEN_1802;
  wire [3:0] _GEN_1803;
  wire [3:0] _GEN_1804;
  wire [3:0] _GEN_1805;
  wire [3:0] _GEN_1806;
  wire [3:0] _GEN_1807;
  wire [3:0] _GEN_1808;
  wire [3:0] _GEN_1809;
  wire [3:0] _GEN_1810;
  wire [3:0] _GEN_1811;
  wire [3:0] _GEN_1812;
  wire [3:0] _GEN_1813;
  wire [3:0] _GEN_1814;
  wire [3:0] _GEN_1815;
  wire [3:0] _GEN_1816;
  wire [3:0] _GEN_1817;
  wire [3:0] _GEN_1818;
  wire [3:0] _GEN_1819;
  wire [3:0] _GEN_1820;
  wire [3:0] _GEN_1821;
  wire [3:0] _GEN_1822;
  wire [3:0] _GEN_1823;
  wire [3:0] _GEN_1824;
  wire [3:0] _GEN_1825;
  wire [6:0] _T_292;
  wire [5:0] _T_293;
  wire [3:0] _T_295;
  wire [3:0] _GEN_28;
  wire [3:0] _GEN_1826;
  wire [3:0] _GEN_1827;
  wire [3:0] _GEN_1828;
  wire [3:0] _GEN_1829;
  wire [3:0] _GEN_1830;
  wire [3:0] _GEN_1831;
  wire [3:0] _GEN_1832;
  wire [3:0] _GEN_1833;
  wire [3:0] _GEN_1834;
  wire [3:0] _GEN_1835;
  wire [3:0] _GEN_1836;
  wire [3:0] _GEN_1837;
  wire [3:0] _GEN_1838;
  wire [3:0] _GEN_1839;
  wire [3:0] _GEN_1840;
  wire [3:0] _GEN_1841;
  wire [3:0] _GEN_1842;
  wire [3:0] _GEN_1843;
  wire [3:0] _GEN_1844;
  wire [3:0] _GEN_1845;
  wire [3:0] _GEN_1846;
  wire [3:0] _GEN_1847;
  wire [3:0] _GEN_1848;
  wire [3:0] _GEN_1849;
  wire [3:0] _GEN_1850;
  wire [3:0] _GEN_1851;
  wire [3:0] _GEN_1852;
  wire [3:0] _GEN_1853;
  wire [3:0] _GEN_1854;
  wire [3:0] _GEN_1855;
  wire [3:0] _GEN_1856;
  wire [3:0] _GEN_1857;
  wire [3:0] _GEN_1858;
  wire [3:0] _GEN_1859;
  wire [3:0] _GEN_1860;
  wire [3:0] _GEN_1861;
  wire [3:0] _GEN_1862;
  wire [3:0] _GEN_1863;
  wire [3:0] _GEN_1864;
  wire [3:0] _GEN_1865;
  wire [3:0] _GEN_1866;
  wire [3:0] _GEN_1867;
  wire [3:0] _GEN_1868;
  wire [3:0] _GEN_1869;
  wire [3:0] _GEN_1870;
  wire [3:0] _GEN_1871;
  wire [3:0] _GEN_1872;
  wire [3:0] _GEN_1873;
  wire [3:0] _GEN_1874;
  wire [3:0] _GEN_1875;
  wire [3:0] _GEN_1876;
  wire [3:0] _GEN_1877;
  wire [3:0] _GEN_1878;
  wire [3:0] _GEN_1879;
  wire [3:0] _GEN_1880;
  wire [3:0] _GEN_1881;
  wire [3:0] _GEN_1882;
  wire [3:0] _GEN_1883;
  wire [3:0] _GEN_1884;
  wire [3:0] _GEN_1885;
  wire [3:0] _GEN_1886;
  wire [3:0] _GEN_1887;
  wire [3:0] _GEN_1888;
  wire [3:0] _GEN_1889;
  wire [6:0] _T_297;
  wire [5:0] _T_298;
  wire [3:0] _T_300;
  wire [3:0] _GEN_29;
  wire [3:0] _GEN_1890;
  wire [3:0] _GEN_1891;
  wire [3:0] _GEN_1892;
  wire [3:0] _GEN_1893;
  wire [3:0] _GEN_1894;
  wire [3:0] _GEN_1895;
  wire [3:0] _GEN_1896;
  wire [3:0] _GEN_1897;
  wire [3:0] _GEN_1898;
  wire [3:0] _GEN_1899;
  wire [3:0] _GEN_1900;
  wire [3:0] _GEN_1901;
  wire [3:0] _GEN_1902;
  wire [3:0] _GEN_1903;
  wire [3:0] _GEN_1904;
  wire [3:0] _GEN_1905;
  wire [3:0] _GEN_1906;
  wire [3:0] _GEN_1907;
  wire [3:0] _GEN_1908;
  wire [3:0] _GEN_1909;
  wire [3:0] _GEN_1910;
  wire [3:0] _GEN_1911;
  wire [3:0] _GEN_1912;
  wire [3:0] _GEN_1913;
  wire [3:0] _GEN_1914;
  wire [3:0] _GEN_1915;
  wire [3:0] _GEN_1916;
  wire [3:0] _GEN_1917;
  wire [3:0] _GEN_1918;
  wire [3:0] _GEN_1919;
  wire [3:0] _GEN_1920;
  wire [3:0] _GEN_1921;
  wire [3:0] _GEN_1922;
  wire [3:0] _GEN_1923;
  wire [3:0] _GEN_1924;
  wire [3:0] _GEN_1925;
  wire [3:0] _GEN_1926;
  wire [3:0] _GEN_1927;
  wire [3:0] _GEN_1928;
  wire [3:0] _GEN_1929;
  wire [3:0] _GEN_1930;
  wire [3:0] _GEN_1931;
  wire [3:0] _GEN_1932;
  wire [3:0] _GEN_1933;
  wire [3:0] _GEN_1934;
  wire [3:0] _GEN_1935;
  wire [3:0] _GEN_1936;
  wire [3:0] _GEN_1937;
  wire [3:0] _GEN_1938;
  wire [3:0] _GEN_1939;
  wire [3:0] _GEN_1940;
  wire [3:0] _GEN_1941;
  wire [3:0] _GEN_1942;
  wire [3:0] _GEN_1943;
  wire [3:0] _GEN_1944;
  wire [3:0] _GEN_1945;
  wire [3:0] _GEN_1946;
  wire [3:0] _GEN_1947;
  wire [3:0] _GEN_1948;
  wire [3:0] _GEN_1949;
  wire [3:0] _GEN_1950;
  wire [3:0] _GEN_1951;
  wire [3:0] _GEN_1952;
  wire [3:0] _GEN_1953;
  wire [6:0] _T_302;
  wire [5:0] _T_303;
  wire [3:0] _T_305;
  wire [3:0] _GEN_30;
  wire [3:0] _GEN_1954;
  wire [3:0] _GEN_1955;
  wire [3:0] _GEN_1956;
  wire [3:0] _GEN_1957;
  wire [3:0] _GEN_1958;
  wire [3:0] _GEN_1959;
  wire [3:0] _GEN_1960;
  wire [3:0] _GEN_1961;
  wire [3:0] _GEN_1962;
  wire [3:0] _GEN_1963;
  wire [3:0] _GEN_1964;
  wire [3:0] _GEN_1965;
  wire [3:0] _GEN_1966;
  wire [3:0] _GEN_1967;
  wire [3:0] _GEN_1968;
  wire [3:0] _GEN_1969;
  wire [3:0] _GEN_1970;
  wire [3:0] _GEN_1971;
  wire [3:0] _GEN_1972;
  wire [3:0] _GEN_1973;
  wire [3:0] _GEN_1974;
  wire [3:0] _GEN_1975;
  wire [3:0] _GEN_1976;
  wire [3:0] _GEN_1977;
  wire [3:0] _GEN_1978;
  wire [3:0] _GEN_1979;
  wire [3:0] _GEN_1980;
  wire [3:0] _GEN_1981;
  wire [3:0] _GEN_1982;
  wire [3:0] _GEN_1983;
  wire [3:0] _GEN_1984;
  wire [3:0] _GEN_1985;
  wire [3:0] _GEN_1986;
  wire [3:0] _GEN_1987;
  wire [3:0] _GEN_1988;
  wire [3:0] _GEN_1989;
  wire [3:0] _GEN_1990;
  wire [3:0] _GEN_1991;
  wire [3:0] _GEN_1992;
  wire [3:0] _GEN_1993;
  wire [3:0] _GEN_1994;
  wire [3:0] _GEN_1995;
  wire [3:0] _GEN_1996;
  wire [3:0] _GEN_1997;
  wire [3:0] _GEN_1998;
  wire [3:0] _GEN_1999;
  wire [3:0] _GEN_2000;
  wire [3:0] _GEN_2001;
  wire [3:0] _GEN_2002;
  wire [3:0] _GEN_2003;
  wire [3:0] _GEN_2004;
  wire [3:0] _GEN_2005;
  wire [3:0] _GEN_2006;
  wire [3:0] _GEN_2007;
  wire [3:0] _GEN_2008;
  wire [3:0] _GEN_2009;
  wire [3:0] _GEN_2010;
  wire [3:0] _GEN_2011;
  wire [3:0] _GEN_2012;
  wire [3:0] _GEN_2013;
  wire [3:0] _GEN_2014;
  wire [3:0] _GEN_2015;
  wire [3:0] _GEN_2016;
  wire [3:0] _GEN_2017;
  wire [6:0] _T_307;
  wire [5:0] _T_308;
  wire [3:0] _T_310;
  wire [3:0] _GEN_31;
  wire [3:0] _GEN_2018;
  wire [3:0] _GEN_2019;
  wire [3:0] _GEN_2020;
  wire [3:0] _GEN_2021;
  wire [3:0] _GEN_2022;
  wire [3:0] _GEN_2023;
  wire [3:0] _GEN_2024;
  wire [3:0] _GEN_2025;
  wire [3:0] _GEN_2026;
  wire [3:0] _GEN_2027;
  wire [3:0] _GEN_2028;
  wire [3:0] _GEN_2029;
  wire [3:0] _GEN_2030;
  wire [3:0] _GEN_2031;
  wire [3:0] _GEN_2032;
  wire [3:0] _GEN_2033;
  wire [3:0] _GEN_2034;
  wire [3:0] _GEN_2035;
  wire [3:0] _GEN_2036;
  wire [3:0] _GEN_2037;
  wire [3:0] _GEN_2038;
  wire [3:0] _GEN_2039;
  wire [3:0] _GEN_2040;
  wire [3:0] _GEN_2041;
  wire [3:0] _GEN_2042;
  wire [3:0] _GEN_2043;
  wire [3:0] _GEN_2044;
  wire [3:0] _GEN_2045;
  wire [3:0] _GEN_2046;
  wire [3:0] _GEN_2047;
  wire [3:0] _GEN_2048;
  wire [3:0] _GEN_2049;
  wire [3:0] _GEN_2050;
  wire [3:0] _GEN_2051;
  wire [3:0] _GEN_2052;
  wire [3:0] _GEN_2053;
  wire [3:0] _GEN_2054;
  wire [3:0] _GEN_2055;
  wire [3:0] _GEN_2056;
  wire [3:0] _GEN_2057;
  wire [3:0] _GEN_2058;
  wire [3:0] _GEN_2059;
  wire [3:0] _GEN_2060;
  wire [3:0] _GEN_2061;
  wire [3:0] _GEN_2062;
  wire [3:0] _GEN_2063;
  wire [3:0] _GEN_2064;
  wire [3:0] _GEN_2065;
  wire [3:0] _GEN_2066;
  wire [3:0] _GEN_2067;
  wire [3:0] _GEN_2068;
  wire [3:0] _GEN_2069;
  wire [3:0] _GEN_2070;
  wire [3:0] _GEN_2071;
  wire [3:0] _GEN_2072;
  wire [3:0] _GEN_2073;
  wire [3:0] _GEN_2074;
  wire [3:0] _GEN_2075;
  wire [3:0] _GEN_2076;
  wire [3:0] _GEN_2077;
  wire [3:0] _GEN_2078;
  wire [3:0] _GEN_2079;
  wire [3:0] _GEN_2080;
  wire [3:0] _GEN_2081;
  wire [6:0] _T_312;
  wire [5:0] _T_313;
  wire [3:0] _GEN_2082;
  wire [3:0] _GEN_2083;
  wire [3:0] _GEN_2084;
  wire [3:0] _GEN_2085;
  wire [3:0] _GEN_2086;
  wire [3:0] _GEN_2087;
  wire [3:0] _GEN_2088;
  wire [3:0] _GEN_2089;
  wire [3:0] _GEN_2090;
  wire [3:0] _GEN_2091;
  wire [3:0] _GEN_2092;
  wire [3:0] _GEN_2093;
  wire [3:0] _GEN_2094;
  wire [3:0] _GEN_2095;
  wire [3:0] _GEN_2096;
  wire [3:0] _GEN_2097;
  wire [3:0] _GEN_2098;
  wire [3:0] _GEN_2099;
  wire [3:0] _GEN_2100;
  wire [3:0] _GEN_2101;
  wire [3:0] _GEN_2102;
  wire [3:0] _GEN_2103;
  wire [3:0] _GEN_2104;
  wire [3:0] _GEN_2105;
  wire [3:0] _GEN_2106;
  wire [3:0] _GEN_2107;
  wire [3:0] _GEN_2108;
  wire [3:0] _GEN_2109;
  wire [3:0] _GEN_2110;
  wire [3:0] _GEN_2111;
  wire [3:0] _GEN_2112;
  wire [3:0] _GEN_2113;
  wire [3:0] _GEN_2114;
  wire [3:0] _GEN_2115;
  wire [3:0] _GEN_2116;
  wire [3:0] _GEN_2117;
  wire [3:0] _GEN_2118;
  wire [3:0] _GEN_2119;
  wire [3:0] _GEN_2120;
  wire [3:0] _GEN_2121;
  wire [3:0] _GEN_2122;
  wire [3:0] _GEN_2123;
  wire [3:0] _GEN_2124;
  wire [3:0] _GEN_2125;
  wire [3:0] _GEN_2126;
  wire [3:0] _GEN_2127;
  wire [3:0] _GEN_2128;
  wire [3:0] _GEN_2129;
  wire [3:0] _GEN_2130;
  wire [3:0] _GEN_2131;
  wire [3:0] _GEN_2132;
  wire [3:0] _GEN_2133;
  wire [3:0] _GEN_2134;
  wire [3:0] _GEN_2135;
  wire [3:0] _GEN_2136;
  wire [3:0] _GEN_2137;
  wire [3:0] _GEN_2138;
  wire [3:0] _GEN_2139;
  wire [3:0] _GEN_2140;
  wire [3:0] _GEN_2141;
  wire [3:0] _GEN_2142;
  wire [3:0] _GEN_2143;
  wire [3:0] _GEN_2144;
  wire [3:0] _GEN_2145;
  wire [5:0] _GEN_2146;
  wire  _T_315;
  wire [3:0] _GEN_32;
  wire [3:0] _GEN_2147;
  wire [3:0] _GEN_2148;
  wire [3:0] _GEN_2149;
  wire [3:0] _GEN_2150;
  wire [3:0] _GEN_2151;
  wire [3:0] _GEN_2152;
  wire [3:0] _GEN_2153;
  wire [3:0] _GEN_2154;
  wire [3:0] _GEN_2155;
  wire [3:0] _GEN_2156;
  wire [3:0] _GEN_2157;
  wire [3:0] _GEN_2158;
  wire [3:0] _GEN_2159;
  wire [3:0] _GEN_2160;
  wire [3:0] _GEN_2161;
  wire [3:0] _GEN_2162;
  wire [3:0] _GEN_2163;
  wire [3:0] _GEN_2164;
  wire [3:0] _GEN_2165;
  wire [3:0] _GEN_2166;
  wire [3:0] _GEN_2167;
  wire [3:0] _GEN_2168;
  wire [3:0] _GEN_2169;
  wire [3:0] _GEN_2170;
  wire [3:0] _GEN_2171;
  wire [3:0] _GEN_2172;
  wire [3:0] _GEN_2173;
  wire [3:0] _GEN_2174;
  wire [3:0] _GEN_2175;
  wire [3:0] _GEN_2176;
  wire [3:0] _GEN_2177;
  wire [3:0] _GEN_2178;
  wire [3:0] _GEN_2179;
  wire [3:0] _GEN_2180;
  wire [3:0] _GEN_2181;
  wire [3:0] _GEN_2182;
  wire [3:0] _GEN_2183;
  wire [3:0] _GEN_2184;
  wire [3:0] _GEN_2185;
  wire [3:0] _GEN_2186;
  wire [3:0] _GEN_2187;
  wire [3:0] _GEN_2188;
  wire [3:0] _GEN_2189;
  wire [3:0] _GEN_2190;
  wire [3:0] _GEN_2191;
  wire [3:0] _GEN_2192;
  wire [3:0] _GEN_2193;
  wire [3:0] _GEN_2194;
  wire [3:0] _GEN_2195;
  wire [3:0] _GEN_2196;
  wire [3:0] _GEN_2197;
  wire [3:0] _GEN_2198;
  wire [3:0] _GEN_2199;
  wire [3:0] _GEN_2200;
  wire [3:0] _GEN_2201;
  wire [3:0] _GEN_2202;
  wire [3:0] _GEN_2203;
  wire [3:0] _GEN_2204;
  wire [3:0] _GEN_2205;
  wire [3:0] _GEN_2206;
  wire [3:0] _GEN_2207;
  wire [3:0] _GEN_2208;
  wire [3:0] _GEN_2209;
  wire [3:0] _GEN_2210;
  wire [3:0] _GEN_2211;
  wire [3:0] _GEN_2212;
  wire [3:0] _GEN_2213;
  wire [3:0] _GEN_2214;
  wire [3:0] _GEN_2215;
  wire [3:0] _GEN_2216;
  wire [3:0] _GEN_2217;
  wire [3:0] _GEN_2218;
  wire [3:0] _GEN_2219;
  wire [3:0] _GEN_2220;
  wire [3:0] _GEN_2221;
  wire [3:0] _GEN_2222;
  wire [3:0] _GEN_2223;
  wire [3:0] _GEN_2224;
  wire [3:0] _GEN_2225;
  wire [3:0] _GEN_2226;
  wire [3:0] _GEN_2227;
  wire [3:0] _GEN_2228;
  wire [3:0] _GEN_2229;
  wire [3:0] _GEN_2230;
  wire [3:0] _GEN_2231;
  wire [3:0] _GEN_2232;
  wire [3:0] _GEN_2233;
  wire [3:0] _GEN_2234;
  wire [3:0] _GEN_2235;
  wire [3:0] _GEN_2236;
  wire [3:0] _GEN_2237;
  wire [3:0] _GEN_2238;
  wire [3:0] _GEN_2239;
  wire [3:0] _GEN_2240;
  wire [3:0] _GEN_2241;
  wire [3:0] _GEN_2242;
  wire [3:0] _GEN_2243;
  wire [3:0] _GEN_2244;
  wire [3:0] _GEN_2245;
  wire [3:0] _GEN_2246;
  wire [3:0] _GEN_2247;
  wire [3:0] _GEN_2248;
  wire [3:0] _GEN_2249;
  wire [3:0] _GEN_2250;
  wire [3:0] _GEN_2251;
  wire [3:0] _GEN_2252;
  wire [3:0] _GEN_2253;
  wire [3:0] _GEN_2254;
  wire [3:0] _GEN_2255;
  wire [3:0] _GEN_2256;
  wire [3:0] _GEN_2257;
  wire [3:0] _GEN_2258;
  wire [3:0] _GEN_2259;
  wire [3:0] _GEN_2260;
  wire [3:0] _GEN_2261;
  wire [3:0] _GEN_2262;
  wire [3:0] _GEN_2263;
  wire [3:0] _GEN_2264;
  wire [3:0] _GEN_2265;
  wire [3:0] _GEN_2266;
  wire [3:0] _GEN_2267;
  wire [3:0] _GEN_2268;
  wire [3:0] _GEN_2269;
  wire [3:0] _GEN_2270;
  wire [3:0] _GEN_2271;
  wire [3:0] _GEN_2272;
  wire [3:0] _GEN_2273;
  wire [3:0] _GEN_2274;
  wire [5:0] _GEN_2275;
  wire  _T_323;
  wire [3:0] _GEN_2276;
  wire [5:0] _GEN_2277;
  wire [2:0] _GEN_2278;
  wire [3:0] _GEN_2279;
  wire [3:0] _GEN_2280;
  wire [3:0] _GEN_2281;
  wire [3:0] _GEN_2282;
  wire [3:0] _GEN_2283;
  wire [3:0] _GEN_2284;
  wire [3:0] _GEN_2285;
  wire [3:0] _GEN_2286;
  wire [3:0] _GEN_2287;
  wire [3:0] _GEN_2288;
  wire [3:0] _GEN_2289;
  wire [3:0] _GEN_2290;
  wire [3:0] _GEN_2291;
  wire [3:0] _GEN_2292;
  wire [3:0] _GEN_2293;
  wire [3:0] _GEN_2294;
  wire [3:0] _GEN_2295;
  wire [3:0] _GEN_2296;
  wire [3:0] _GEN_2297;
  wire [3:0] _GEN_2298;
  wire [3:0] _GEN_2299;
  wire [3:0] _GEN_2300;
  wire [3:0] _GEN_2301;
  wire [3:0] _GEN_2302;
  wire [3:0] _GEN_2303;
  wire [3:0] _GEN_2304;
  wire [3:0] _GEN_2305;
  wire [3:0] _GEN_2306;
  wire [3:0] _GEN_2307;
  wire [3:0] _GEN_2308;
  wire [3:0] _GEN_2309;
  wire [3:0] _GEN_2310;
  wire [3:0] _GEN_2311;
  wire [3:0] _GEN_2312;
  wire [3:0] _GEN_2313;
  wire [3:0] _GEN_2314;
  wire [3:0] _GEN_2315;
  wire [3:0] _GEN_2316;
  wire [3:0] _GEN_2317;
  wire [3:0] _GEN_2318;
  wire [3:0] _GEN_2319;
  wire [3:0] _GEN_2320;
  wire [3:0] _GEN_2321;
  wire [3:0] _GEN_2322;
  wire [3:0] _GEN_2323;
  wire [3:0] _GEN_2324;
  wire [3:0] _GEN_2325;
  wire [3:0] _GEN_2326;
  wire [3:0] _GEN_2327;
  wire [3:0] _GEN_2328;
  wire [3:0] _GEN_2329;
  wire [3:0] _GEN_2330;
  wire [3:0] _GEN_2331;
  wire [3:0] _GEN_2332;
  wire [3:0] _GEN_2333;
  wire [3:0] _GEN_2334;
  wire [3:0] _GEN_2335;
  wire [3:0] _GEN_2336;
  wire [3:0] _GEN_2337;
  wire [3:0] _GEN_2338;
  wire [3:0] _GEN_2339;
  wire [3:0] _GEN_2340;
  wire [3:0] _GEN_2341;
  wire [3:0] _GEN_2342;
  wire [5:0] _GEN_2343;
  wire [2:0] _GEN_2344;
  wire [3:0] _T_329;
  wire [2:0] _T_330;
  wire [2:0] _GEN_2345;
  wire [2:0] _GEN_2346;
  wire [5:0] _GEN_2347;
  wire [2:0] _GEN_2348;
  wire [5:0] _GEN_2349;
  wire [3:0] _GEN_2350;
  wire [3:0] _GEN_2351;
  wire [3:0] _GEN_2352;
  wire [3:0] _GEN_2353;
  wire [3:0] _GEN_2354;
  wire [3:0] _GEN_2355;
  wire [3:0] _GEN_2356;
  wire [3:0] _GEN_2357;
  wire [3:0] _GEN_2358;
  wire [3:0] _GEN_2359;
  wire [3:0] _GEN_2360;
  wire [3:0] _GEN_2361;
  wire [3:0] _GEN_2362;
  wire [3:0] _GEN_2363;
  wire [3:0] _GEN_2364;
  wire [3:0] _GEN_2365;
  wire [3:0] _GEN_2366;
  wire [3:0] _GEN_2367;
  wire [3:0] _GEN_2368;
  wire [3:0] _GEN_2369;
  wire [3:0] _GEN_2370;
  wire [3:0] _GEN_2371;
  wire [3:0] _GEN_2372;
  wire [3:0] _GEN_2373;
  wire [3:0] _GEN_2374;
  wire [3:0] _GEN_2375;
  wire [3:0] _GEN_2376;
  wire [3:0] _GEN_2377;
  wire [3:0] _GEN_2378;
  wire [3:0] _GEN_2379;
  wire [3:0] _GEN_2380;
  wire [3:0] _GEN_2381;
  wire [3:0] _GEN_2382;
  wire [3:0] _GEN_2383;
  wire [3:0] _GEN_2384;
  wire [3:0] _GEN_2385;
  wire [3:0] _GEN_2386;
  wire [3:0] _GEN_2387;
  wire [3:0] _GEN_2388;
  wire [3:0] _GEN_2389;
  wire [3:0] _GEN_2390;
  wire [3:0] _GEN_2391;
  wire [3:0] _GEN_2392;
  wire [3:0] _GEN_2393;
  wire [3:0] _GEN_2394;
  wire [3:0] _GEN_2395;
  wire [3:0] _GEN_2396;
  wire [3:0] _GEN_2397;
  wire [3:0] _GEN_2398;
  wire [3:0] _GEN_2399;
  wire [3:0] _GEN_2400;
  wire [3:0] _GEN_2401;
  wire [3:0] _GEN_2402;
  wire [3:0] _GEN_2403;
  wire [3:0] _GEN_2404;
  wire [3:0] _GEN_2405;
  wire [3:0] _GEN_2406;
  wire [3:0] _GEN_2407;
  wire [3:0] _GEN_2408;
  wire [3:0] _GEN_2409;
  wire [3:0] _GEN_2410;
  wire [3:0] _GEN_2411;
  wire [3:0] _GEN_2412;
  wire [3:0] _GEN_2413;
  wire [5:0] _GEN_2414;
  wire [2:0] _GEN_2415;
  wire  _T_336;
  wire  _T_337;
  wire  _T_339;
  wire  _T_340;
  wire [5:0] _GEN_2416;
  wire [2:0] _GEN_2417;
  wire [31:0] _GEN_33;
  wire [31:0] _GEN_2418;
  wire [31:0] _GEN_2419;
  wire [31:0] _GEN_2420;
  wire [31:0] _GEN_2421;
  wire [31:0] _GEN_2422;
  wire [31:0] _GEN_2423;
  wire [31:0] _GEN_2424;
  assign io_out = _GEN_33;
  assign _T_80 = {mem_6,mem_7};
  assign _T_81 = {mem_4,mem_5};
  assign _T_82 = {_T_81,_T_80};
  assign _T_83 = {mem_2,mem_3};
  assign _T_84 = {mem_0,mem_1};
  assign _T_85 = {_T_84,_T_83};
  assign _T_86 = {_T_85,_T_82};
  assign _T_87 = {mem_14,mem_15};
  assign _T_88 = {mem_12,mem_13};
  assign _T_89 = {_T_88,_T_87};
  assign _T_90 = {mem_10,mem_11};
  assign _T_91 = {mem_8,mem_9};
  assign _T_92 = {_T_91,_T_90};
  assign _T_93 = {_T_92,_T_89};
  assign _T_94 = {mem_22,mem_23};
  assign _T_95 = {mem_20,mem_21};
  assign _T_96 = {_T_95,_T_94};
  assign _T_97 = {mem_18,mem_19};
  assign _T_98 = {mem_16,mem_17};
  assign _T_99 = {_T_98,_T_97};
  assign _T_100 = {_T_99,_T_96};
  assign _T_101 = {mem_30,mem_31};
  assign _T_102 = {mem_28,mem_29};
  assign _T_103 = {_T_102,_T_101};
  assign _T_104 = {mem_26,mem_27};
  assign _T_105 = {mem_24,mem_25};
  assign _T_106 = {_T_105,_T_104};
  assign _T_107 = {_T_106,_T_103};
  assign _T_108 = {mem_38,mem_39};
  assign _T_109 = {mem_36,mem_37};
  assign _T_110 = {_T_109,_T_108};
  assign _T_111 = {mem_34,mem_35};
  assign _T_112 = {mem_32,mem_33};
  assign _T_113 = {_T_112,_T_111};
  assign _T_114 = {_T_113,_T_110};
  assign _T_115 = {mem_46,mem_47};
  assign _T_116 = {mem_44,mem_45};
  assign _T_117 = {_T_116,_T_115};
  assign _T_118 = {mem_42,mem_43};
  assign _T_119 = {mem_40,mem_41};
  assign _T_120 = {_T_119,_T_118};
  assign _T_121 = {_T_120,_T_117};
  assign _T_122 = {mem_54,mem_55};
  assign _T_123 = {mem_52,mem_53};
  assign _T_124 = {_T_123,_T_122};
  assign _T_125 = {mem_50,mem_51};
  assign _T_126 = {mem_48,mem_49};
  assign _T_127 = {_T_126,_T_125};
  assign _T_128 = {_T_127,_T_124};
  assign _T_129 = {mem_62,mem_63};
  assign _T_130 = {mem_60,mem_61};
  assign _T_131 = {_T_130,_T_129};
  assign _T_132 = {mem_58,mem_59};
  assign _T_133 = {mem_56,mem_57};
  assign _T_134 = {_T_133,_T_132};
  assign _T_135 = {_T_134,_T_131};
  assign catMem_0 = _T_86;
  assign catMem_1 = _T_93;
  assign catMem_2 = _T_100;
  assign catMem_3 = _T_107;
  assign catMem_4 = _T_114;
  assign catMem_5 = _T_121;
  assign catMem_6 = _T_128;
  assign catMem_7 = _T_135;
  assign _T_149 = io_reset == 1'h0;
  assign _T_150 = io_fastpush & _T_149;
  assign _T_152 = wPos + 6'h0;
  assign _T_153 = _T_152[5:0];
  assign _T_155 = io_fastin[127:124];
  assign _GEN_0 = _T_155;
  assign _GEN_34 = 6'h0 == _T_153 ? _GEN_0 : mem_0;
  assign _GEN_35 = 6'h1 == _T_153 ? _GEN_0 : mem_1;
  assign _GEN_36 = 6'h2 == _T_153 ? _GEN_0 : mem_2;
  assign _GEN_37 = 6'h3 == _T_153 ? _GEN_0 : mem_3;
  assign _GEN_38 = 6'h4 == _T_153 ? _GEN_0 : mem_4;
  assign _GEN_39 = 6'h5 == _T_153 ? _GEN_0 : mem_5;
  assign _GEN_40 = 6'h6 == _T_153 ? _GEN_0 : mem_6;
  assign _GEN_41 = 6'h7 == _T_153 ? _GEN_0 : mem_7;
  assign _GEN_42 = 6'h8 == _T_153 ? _GEN_0 : mem_8;
  assign _GEN_43 = 6'h9 == _T_153 ? _GEN_0 : mem_9;
  assign _GEN_44 = 6'ha == _T_153 ? _GEN_0 : mem_10;
  assign _GEN_45 = 6'hb == _T_153 ? _GEN_0 : mem_11;
  assign _GEN_46 = 6'hc == _T_153 ? _GEN_0 : mem_12;
  assign _GEN_47 = 6'hd == _T_153 ? _GEN_0 : mem_13;
  assign _GEN_48 = 6'he == _T_153 ? _GEN_0 : mem_14;
  assign _GEN_49 = 6'hf == _T_153 ? _GEN_0 : mem_15;
  assign _GEN_50 = 6'h10 == _T_153 ? _GEN_0 : mem_16;
  assign _GEN_51 = 6'h11 == _T_153 ? _GEN_0 : mem_17;
  assign _GEN_52 = 6'h12 == _T_153 ? _GEN_0 : mem_18;
  assign _GEN_53 = 6'h13 == _T_153 ? _GEN_0 : mem_19;
  assign _GEN_54 = 6'h14 == _T_153 ? _GEN_0 : mem_20;
  assign _GEN_55 = 6'h15 == _T_153 ? _GEN_0 : mem_21;
  assign _GEN_56 = 6'h16 == _T_153 ? _GEN_0 : mem_22;
  assign _GEN_57 = 6'h17 == _T_153 ? _GEN_0 : mem_23;
  assign _GEN_58 = 6'h18 == _T_153 ? _GEN_0 : mem_24;
  assign _GEN_59 = 6'h19 == _T_153 ? _GEN_0 : mem_25;
  assign _GEN_60 = 6'h1a == _T_153 ? _GEN_0 : mem_26;
  assign _GEN_61 = 6'h1b == _T_153 ? _GEN_0 : mem_27;
  assign _GEN_62 = 6'h1c == _T_153 ? _GEN_0 : mem_28;
  assign _GEN_63 = 6'h1d == _T_153 ? _GEN_0 : mem_29;
  assign _GEN_64 = 6'h1e == _T_153 ? _GEN_0 : mem_30;
  assign _GEN_65 = 6'h1f == _T_153 ? _GEN_0 : mem_31;
  assign _GEN_66 = 6'h20 == _T_153 ? _GEN_0 : mem_32;
  assign _GEN_67 = 6'h21 == _T_153 ? _GEN_0 : mem_33;
  assign _GEN_68 = 6'h22 == _T_153 ? _GEN_0 : mem_34;
  assign _GEN_69 = 6'h23 == _T_153 ? _GEN_0 : mem_35;
  assign _GEN_70 = 6'h24 == _T_153 ? _GEN_0 : mem_36;
  assign _GEN_71 = 6'h25 == _T_153 ? _GEN_0 : mem_37;
  assign _GEN_72 = 6'h26 == _T_153 ? _GEN_0 : mem_38;
  assign _GEN_73 = 6'h27 == _T_153 ? _GEN_0 : mem_39;
  assign _GEN_74 = 6'h28 == _T_153 ? _GEN_0 : mem_40;
  assign _GEN_75 = 6'h29 == _T_153 ? _GEN_0 : mem_41;
  assign _GEN_76 = 6'h2a == _T_153 ? _GEN_0 : mem_42;
  assign _GEN_77 = 6'h2b == _T_153 ? _GEN_0 : mem_43;
  assign _GEN_78 = 6'h2c == _T_153 ? _GEN_0 : mem_44;
  assign _GEN_79 = 6'h2d == _T_153 ? _GEN_0 : mem_45;
  assign _GEN_80 = 6'h2e == _T_153 ? _GEN_0 : mem_46;
  assign _GEN_81 = 6'h2f == _T_153 ? _GEN_0 : mem_47;
  assign _GEN_82 = 6'h30 == _T_153 ? _GEN_0 : mem_48;
  assign _GEN_83 = 6'h31 == _T_153 ? _GEN_0 : mem_49;
  assign _GEN_84 = 6'h32 == _T_153 ? _GEN_0 : mem_50;
  assign _GEN_85 = 6'h33 == _T_153 ? _GEN_0 : mem_51;
  assign _GEN_86 = 6'h34 == _T_153 ? _GEN_0 : mem_52;
  assign _GEN_87 = 6'h35 == _T_153 ? _GEN_0 : mem_53;
  assign _GEN_88 = 6'h36 == _T_153 ? _GEN_0 : mem_54;
  assign _GEN_89 = 6'h37 == _T_153 ? _GEN_0 : mem_55;
  assign _GEN_90 = 6'h38 == _T_153 ? _GEN_0 : mem_56;
  assign _GEN_91 = 6'h39 == _T_153 ? _GEN_0 : mem_57;
  assign _GEN_92 = 6'h3a == _T_153 ? _GEN_0 : mem_58;
  assign _GEN_93 = 6'h3b == _T_153 ? _GEN_0 : mem_59;
  assign _GEN_94 = 6'h3c == _T_153 ? _GEN_0 : mem_60;
  assign _GEN_95 = 6'h3d == _T_153 ? _GEN_0 : mem_61;
  assign _GEN_96 = 6'h3e == _T_153 ? _GEN_0 : mem_62;
  assign _GEN_97 = 6'h3f == _T_153 ? _GEN_0 : mem_63;
  assign _T_157 = wPos + 6'h1;
  assign _T_158 = _T_157[5:0];
  assign _T_160 = io_fastin[123:120];
  assign _GEN_1 = _T_160;
  assign _GEN_98 = 6'h0 == _T_158 ? _GEN_1 : _GEN_34;
  assign _GEN_99 = 6'h1 == _T_158 ? _GEN_1 : _GEN_35;
  assign _GEN_100 = 6'h2 == _T_158 ? _GEN_1 : _GEN_36;
  assign _GEN_101 = 6'h3 == _T_158 ? _GEN_1 : _GEN_37;
  assign _GEN_102 = 6'h4 == _T_158 ? _GEN_1 : _GEN_38;
  assign _GEN_103 = 6'h5 == _T_158 ? _GEN_1 : _GEN_39;
  assign _GEN_104 = 6'h6 == _T_158 ? _GEN_1 : _GEN_40;
  assign _GEN_105 = 6'h7 == _T_158 ? _GEN_1 : _GEN_41;
  assign _GEN_106 = 6'h8 == _T_158 ? _GEN_1 : _GEN_42;
  assign _GEN_107 = 6'h9 == _T_158 ? _GEN_1 : _GEN_43;
  assign _GEN_108 = 6'ha == _T_158 ? _GEN_1 : _GEN_44;
  assign _GEN_109 = 6'hb == _T_158 ? _GEN_1 : _GEN_45;
  assign _GEN_110 = 6'hc == _T_158 ? _GEN_1 : _GEN_46;
  assign _GEN_111 = 6'hd == _T_158 ? _GEN_1 : _GEN_47;
  assign _GEN_112 = 6'he == _T_158 ? _GEN_1 : _GEN_48;
  assign _GEN_113 = 6'hf == _T_158 ? _GEN_1 : _GEN_49;
  assign _GEN_114 = 6'h10 == _T_158 ? _GEN_1 : _GEN_50;
  assign _GEN_115 = 6'h11 == _T_158 ? _GEN_1 : _GEN_51;
  assign _GEN_116 = 6'h12 == _T_158 ? _GEN_1 : _GEN_52;
  assign _GEN_117 = 6'h13 == _T_158 ? _GEN_1 : _GEN_53;
  assign _GEN_118 = 6'h14 == _T_158 ? _GEN_1 : _GEN_54;
  assign _GEN_119 = 6'h15 == _T_158 ? _GEN_1 : _GEN_55;
  assign _GEN_120 = 6'h16 == _T_158 ? _GEN_1 : _GEN_56;
  assign _GEN_121 = 6'h17 == _T_158 ? _GEN_1 : _GEN_57;
  assign _GEN_122 = 6'h18 == _T_158 ? _GEN_1 : _GEN_58;
  assign _GEN_123 = 6'h19 == _T_158 ? _GEN_1 : _GEN_59;
  assign _GEN_124 = 6'h1a == _T_158 ? _GEN_1 : _GEN_60;
  assign _GEN_125 = 6'h1b == _T_158 ? _GEN_1 : _GEN_61;
  assign _GEN_126 = 6'h1c == _T_158 ? _GEN_1 : _GEN_62;
  assign _GEN_127 = 6'h1d == _T_158 ? _GEN_1 : _GEN_63;
  assign _GEN_128 = 6'h1e == _T_158 ? _GEN_1 : _GEN_64;
  assign _GEN_129 = 6'h1f == _T_158 ? _GEN_1 : _GEN_65;
  assign _GEN_130 = 6'h20 == _T_158 ? _GEN_1 : _GEN_66;
  assign _GEN_131 = 6'h21 == _T_158 ? _GEN_1 : _GEN_67;
  assign _GEN_132 = 6'h22 == _T_158 ? _GEN_1 : _GEN_68;
  assign _GEN_133 = 6'h23 == _T_158 ? _GEN_1 : _GEN_69;
  assign _GEN_134 = 6'h24 == _T_158 ? _GEN_1 : _GEN_70;
  assign _GEN_135 = 6'h25 == _T_158 ? _GEN_1 : _GEN_71;
  assign _GEN_136 = 6'h26 == _T_158 ? _GEN_1 : _GEN_72;
  assign _GEN_137 = 6'h27 == _T_158 ? _GEN_1 : _GEN_73;
  assign _GEN_138 = 6'h28 == _T_158 ? _GEN_1 : _GEN_74;
  assign _GEN_139 = 6'h29 == _T_158 ? _GEN_1 : _GEN_75;
  assign _GEN_140 = 6'h2a == _T_158 ? _GEN_1 : _GEN_76;
  assign _GEN_141 = 6'h2b == _T_158 ? _GEN_1 : _GEN_77;
  assign _GEN_142 = 6'h2c == _T_158 ? _GEN_1 : _GEN_78;
  assign _GEN_143 = 6'h2d == _T_158 ? _GEN_1 : _GEN_79;
  assign _GEN_144 = 6'h2e == _T_158 ? _GEN_1 : _GEN_80;
  assign _GEN_145 = 6'h2f == _T_158 ? _GEN_1 : _GEN_81;
  assign _GEN_146 = 6'h30 == _T_158 ? _GEN_1 : _GEN_82;
  assign _GEN_147 = 6'h31 == _T_158 ? _GEN_1 : _GEN_83;
  assign _GEN_148 = 6'h32 == _T_158 ? _GEN_1 : _GEN_84;
  assign _GEN_149 = 6'h33 == _T_158 ? _GEN_1 : _GEN_85;
  assign _GEN_150 = 6'h34 == _T_158 ? _GEN_1 : _GEN_86;
  assign _GEN_151 = 6'h35 == _T_158 ? _GEN_1 : _GEN_87;
  assign _GEN_152 = 6'h36 == _T_158 ? _GEN_1 : _GEN_88;
  assign _GEN_153 = 6'h37 == _T_158 ? _GEN_1 : _GEN_89;
  assign _GEN_154 = 6'h38 == _T_158 ? _GEN_1 : _GEN_90;
  assign _GEN_155 = 6'h39 == _T_158 ? _GEN_1 : _GEN_91;
  assign _GEN_156 = 6'h3a == _T_158 ? _GEN_1 : _GEN_92;
  assign _GEN_157 = 6'h3b == _T_158 ? _GEN_1 : _GEN_93;
  assign _GEN_158 = 6'h3c == _T_158 ? _GEN_1 : _GEN_94;
  assign _GEN_159 = 6'h3d == _T_158 ? _GEN_1 : _GEN_95;
  assign _GEN_160 = 6'h3e == _T_158 ? _GEN_1 : _GEN_96;
  assign _GEN_161 = 6'h3f == _T_158 ? _GEN_1 : _GEN_97;
  assign _T_162 = wPos + 6'h2;
  assign _T_163 = _T_162[5:0];
  assign _T_165 = io_fastin[119:116];
  assign _GEN_2 = _T_165;
  assign _GEN_162 = 6'h0 == _T_163 ? _GEN_2 : _GEN_98;
  assign _GEN_163 = 6'h1 == _T_163 ? _GEN_2 : _GEN_99;
  assign _GEN_164 = 6'h2 == _T_163 ? _GEN_2 : _GEN_100;
  assign _GEN_165 = 6'h3 == _T_163 ? _GEN_2 : _GEN_101;
  assign _GEN_166 = 6'h4 == _T_163 ? _GEN_2 : _GEN_102;
  assign _GEN_167 = 6'h5 == _T_163 ? _GEN_2 : _GEN_103;
  assign _GEN_168 = 6'h6 == _T_163 ? _GEN_2 : _GEN_104;
  assign _GEN_169 = 6'h7 == _T_163 ? _GEN_2 : _GEN_105;
  assign _GEN_170 = 6'h8 == _T_163 ? _GEN_2 : _GEN_106;
  assign _GEN_171 = 6'h9 == _T_163 ? _GEN_2 : _GEN_107;
  assign _GEN_172 = 6'ha == _T_163 ? _GEN_2 : _GEN_108;
  assign _GEN_173 = 6'hb == _T_163 ? _GEN_2 : _GEN_109;
  assign _GEN_174 = 6'hc == _T_163 ? _GEN_2 : _GEN_110;
  assign _GEN_175 = 6'hd == _T_163 ? _GEN_2 : _GEN_111;
  assign _GEN_176 = 6'he == _T_163 ? _GEN_2 : _GEN_112;
  assign _GEN_177 = 6'hf == _T_163 ? _GEN_2 : _GEN_113;
  assign _GEN_178 = 6'h10 == _T_163 ? _GEN_2 : _GEN_114;
  assign _GEN_179 = 6'h11 == _T_163 ? _GEN_2 : _GEN_115;
  assign _GEN_180 = 6'h12 == _T_163 ? _GEN_2 : _GEN_116;
  assign _GEN_181 = 6'h13 == _T_163 ? _GEN_2 : _GEN_117;
  assign _GEN_182 = 6'h14 == _T_163 ? _GEN_2 : _GEN_118;
  assign _GEN_183 = 6'h15 == _T_163 ? _GEN_2 : _GEN_119;
  assign _GEN_184 = 6'h16 == _T_163 ? _GEN_2 : _GEN_120;
  assign _GEN_185 = 6'h17 == _T_163 ? _GEN_2 : _GEN_121;
  assign _GEN_186 = 6'h18 == _T_163 ? _GEN_2 : _GEN_122;
  assign _GEN_187 = 6'h19 == _T_163 ? _GEN_2 : _GEN_123;
  assign _GEN_188 = 6'h1a == _T_163 ? _GEN_2 : _GEN_124;
  assign _GEN_189 = 6'h1b == _T_163 ? _GEN_2 : _GEN_125;
  assign _GEN_190 = 6'h1c == _T_163 ? _GEN_2 : _GEN_126;
  assign _GEN_191 = 6'h1d == _T_163 ? _GEN_2 : _GEN_127;
  assign _GEN_192 = 6'h1e == _T_163 ? _GEN_2 : _GEN_128;
  assign _GEN_193 = 6'h1f == _T_163 ? _GEN_2 : _GEN_129;
  assign _GEN_194 = 6'h20 == _T_163 ? _GEN_2 : _GEN_130;
  assign _GEN_195 = 6'h21 == _T_163 ? _GEN_2 : _GEN_131;
  assign _GEN_196 = 6'h22 == _T_163 ? _GEN_2 : _GEN_132;
  assign _GEN_197 = 6'h23 == _T_163 ? _GEN_2 : _GEN_133;
  assign _GEN_198 = 6'h24 == _T_163 ? _GEN_2 : _GEN_134;
  assign _GEN_199 = 6'h25 == _T_163 ? _GEN_2 : _GEN_135;
  assign _GEN_200 = 6'h26 == _T_163 ? _GEN_2 : _GEN_136;
  assign _GEN_201 = 6'h27 == _T_163 ? _GEN_2 : _GEN_137;
  assign _GEN_202 = 6'h28 == _T_163 ? _GEN_2 : _GEN_138;
  assign _GEN_203 = 6'h29 == _T_163 ? _GEN_2 : _GEN_139;
  assign _GEN_204 = 6'h2a == _T_163 ? _GEN_2 : _GEN_140;
  assign _GEN_205 = 6'h2b == _T_163 ? _GEN_2 : _GEN_141;
  assign _GEN_206 = 6'h2c == _T_163 ? _GEN_2 : _GEN_142;
  assign _GEN_207 = 6'h2d == _T_163 ? _GEN_2 : _GEN_143;
  assign _GEN_208 = 6'h2e == _T_163 ? _GEN_2 : _GEN_144;
  assign _GEN_209 = 6'h2f == _T_163 ? _GEN_2 : _GEN_145;
  assign _GEN_210 = 6'h30 == _T_163 ? _GEN_2 : _GEN_146;
  assign _GEN_211 = 6'h31 == _T_163 ? _GEN_2 : _GEN_147;
  assign _GEN_212 = 6'h32 == _T_163 ? _GEN_2 : _GEN_148;
  assign _GEN_213 = 6'h33 == _T_163 ? _GEN_2 : _GEN_149;
  assign _GEN_214 = 6'h34 == _T_163 ? _GEN_2 : _GEN_150;
  assign _GEN_215 = 6'h35 == _T_163 ? _GEN_2 : _GEN_151;
  assign _GEN_216 = 6'h36 == _T_163 ? _GEN_2 : _GEN_152;
  assign _GEN_217 = 6'h37 == _T_163 ? _GEN_2 : _GEN_153;
  assign _GEN_218 = 6'h38 == _T_163 ? _GEN_2 : _GEN_154;
  assign _GEN_219 = 6'h39 == _T_163 ? _GEN_2 : _GEN_155;
  assign _GEN_220 = 6'h3a == _T_163 ? _GEN_2 : _GEN_156;
  assign _GEN_221 = 6'h3b == _T_163 ? _GEN_2 : _GEN_157;
  assign _GEN_222 = 6'h3c == _T_163 ? _GEN_2 : _GEN_158;
  assign _GEN_223 = 6'h3d == _T_163 ? _GEN_2 : _GEN_159;
  assign _GEN_224 = 6'h3e == _T_163 ? _GEN_2 : _GEN_160;
  assign _GEN_225 = 6'h3f == _T_163 ? _GEN_2 : _GEN_161;
  assign _T_167 = wPos + 6'h3;
  assign _T_168 = _T_167[5:0];
  assign _T_170 = io_fastin[115:112];
  assign _GEN_3 = _T_170;
  assign _GEN_226 = 6'h0 == _T_168 ? _GEN_3 : _GEN_162;
  assign _GEN_227 = 6'h1 == _T_168 ? _GEN_3 : _GEN_163;
  assign _GEN_228 = 6'h2 == _T_168 ? _GEN_3 : _GEN_164;
  assign _GEN_229 = 6'h3 == _T_168 ? _GEN_3 : _GEN_165;
  assign _GEN_230 = 6'h4 == _T_168 ? _GEN_3 : _GEN_166;
  assign _GEN_231 = 6'h5 == _T_168 ? _GEN_3 : _GEN_167;
  assign _GEN_232 = 6'h6 == _T_168 ? _GEN_3 : _GEN_168;
  assign _GEN_233 = 6'h7 == _T_168 ? _GEN_3 : _GEN_169;
  assign _GEN_234 = 6'h8 == _T_168 ? _GEN_3 : _GEN_170;
  assign _GEN_235 = 6'h9 == _T_168 ? _GEN_3 : _GEN_171;
  assign _GEN_236 = 6'ha == _T_168 ? _GEN_3 : _GEN_172;
  assign _GEN_237 = 6'hb == _T_168 ? _GEN_3 : _GEN_173;
  assign _GEN_238 = 6'hc == _T_168 ? _GEN_3 : _GEN_174;
  assign _GEN_239 = 6'hd == _T_168 ? _GEN_3 : _GEN_175;
  assign _GEN_240 = 6'he == _T_168 ? _GEN_3 : _GEN_176;
  assign _GEN_241 = 6'hf == _T_168 ? _GEN_3 : _GEN_177;
  assign _GEN_242 = 6'h10 == _T_168 ? _GEN_3 : _GEN_178;
  assign _GEN_243 = 6'h11 == _T_168 ? _GEN_3 : _GEN_179;
  assign _GEN_244 = 6'h12 == _T_168 ? _GEN_3 : _GEN_180;
  assign _GEN_245 = 6'h13 == _T_168 ? _GEN_3 : _GEN_181;
  assign _GEN_246 = 6'h14 == _T_168 ? _GEN_3 : _GEN_182;
  assign _GEN_247 = 6'h15 == _T_168 ? _GEN_3 : _GEN_183;
  assign _GEN_248 = 6'h16 == _T_168 ? _GEN_3 : _GEN_184;
  assign _GEN_249 = 6'h17 == _T_168 ? _GEN_3 : _GEN_185;
  assign _GEN_250 = 6'h18 == _T_168 ? _GEN_3 : _GEN_186;
  assign _GEN_251 = 6'h19 == _T_168 ? _GEN_3 : _GEN_187;
  assign _GEN_252 = 6'h1a == _T_168 ? _GEN_3 : _GEN_188;
  assign _GEN_253 = 6'h1b == _T_168 ? _GEN_3 : _GEN_189;
  assign _GEN_254 = 6'h1c == _T_168 ? _GEN_3 : _GEN_190;
  assign _GEN_255 = 6'h1d == _T_168 ? _GEN_3 : _GEN_191;
  assign _GEN_256 = 6'h1e == _T_168 ? _GEN_3 : _GEN_192;
  assign _GEN_257 = 6'h1f == _T_168 ? _GEN_3 : _GEN_193;
  assign _GEN_258 = 6'h20 == _T_168 ? _GEN_3 : _GEN_194;
  assign _GEN_259 = 6'h21 == _T_168 ? _GEN_3 : _GEN_195;
  assign _GEN_260 = 6'h22 == _T_168 ? _GEN_3 : _GEN_196;
  assign _GEN_261 = 6'h23 == _T_168 ? _GEN_3 : _GEN_197;
  assign _GEN_262 = 6'h24 == _T_168 ? _GEN_3 : _GEN_198;
  assign _GEN_263 = 6'h25 == _T_168 ? _GEN_3 : _GEN_199;
  assign _GEN_264 = 6'h26 == _T_168 ? _GEN_3 : _GEN_200;
  assign _GEN_265 = 6'h27 == _T_168 ? _GEN_3 : _GEN_201;
  assign _GEN_266 = 6'h28 == _T_168 ? _GEN_3 : _GEN_202;
  assign _GEN_267 = 6'h29 == _T_168 ? _GEN_3 : _GEN_203;
  assign _GEN_268 = 6'h2a == _T_168 ? _GEN_3 : _GEN_204;
  assign _GEN_269 = 6'h2b == _T_168 ? _GEN_3 : _GEN_205;
  assign _GEN_270 = 6'h2c == _T_168 ? _GEN_3 : _GEN_206;
  assign _GEN_271 = 6'h2d == _T_168 ? _GEN_3 : _GEN_207;
  assign _GEN_272 = 6'h2e == _T_168 ? _GEN_3 : _GEN_208;
  assign _GEN_273 = 6'h2f == _T_168 ? _GEN_3 : _GEN_209;
  assign _GEN_274 = 6'h30 == _T_168 ? _GEN_3 : _GEN_210;
  assign _GEN_275 = 6'h31 == _T_168 ? _GEN_3 : _GEN_211;
  assign _GEN_276 = 6'h32 == _T_168 ? _GEN_3 : _GEN_212;
  assign _GEN_277 = 6'h33 == _T_168 ? _GEN_3 : _GEN_213;
  assign _GEN_278 = 6'h34 == _T_168 ? _GEN_3 : _GEN_214;
  assign _GEN_279 = 6'h35 == _T_168 ? _GEN_3 : _GEN_215;
  assign _GEN_280 = 6'h36 == _T_168 ? _GEN_3 : _GEN_216;
  assign _GEN_281 = 6'h37 == _T_168 ? _GEN_3 : _GEN_217;
  assign _GEN_282 = 6'h38 == _T_168 ? _GEN_3 : _GEN_218;
  assign _GEN_283 = 6'h39 == _T_168 ? _GEN_3 : _GEN_219;
  assign _GEN_284 = 6'h3a == _T_168 ? _GEN_3 : _GEN_220;
  assign _GEN_285 = 6'h3b == _T_168 ? _GEN_3 : _GEN_221;
  assign _GEN_286 = 6'h3c == _T_168 ? _GEN_3 : _GEN_222;
  assign _GEN_287 = 6'h3d == _T_168 ? _GEN_3 : _GEN_223;
  assign _GEN_288 = 6'h3e == _T_168 ? _GEN_3 : _GEN_224;
  assign _GEN_289 = 6'h3f == _T_168 ? _GEN_3 : _GEN_225;
  assign _T_172 = wPos + 6'h4;
  assign _T_173 = _T_172[5:0];
  assign _T_175 = io_fastin[111:108];
  assign _GEN_4 = _T_175;
  assign _GEN_290 = 6'h0 == _T_173 ? _GEN_4 : _GEN_226;
  assign _GEN_291 = 6'h1 == _T_173 ? _GEN_4 : _GEN_227;
  assign _GEN_292 = 6'h2 == _T_173 ? _GEN_4 : _GEN_228;
  assign _GEN_293 = 6'h3 == _T_173 ? _GEN_4 : _GEN_229;
  assign _GEN_294 = 6'h4 == _T_173 ? _GEN_4 : _GEN_230;
  assign _GEN_295 = 6'h5 == _T_173 ? _GEN_4 : _GEN_231;
  assign _GEN_296 = 6'h6 == _T_173 ? _GEN_4 : _GEN_232;
  assign _GEN_297 = 6'h7 == _T_173 ? _GEN_4 : _GEN_233;
  assign _GEN_298 = 6'h8 == _T_173 ? _GEN_4 : _GEN_234;
  assign _GEN_299 = 6'h9 == _T_173 ? _GEN_4 : _GEN_235;
  assign _GEN_300 = 6'ha == _T_173 ? _GEN_4 : _GEN_236;
  assign _GEN_301 = 6'hb == _T_173 ? _GEN_4 : _GEN_237;
  assign _GEN_302 = 6'hc == _T_173 ? _GEN_4 : _GEN_238;
  assign _GEN_303 = 6'hd == _T_173 ? _GEN_4 : _GEN_239;
  assign _GEN_304 = 6'he == _T_173 ? _GEN_4 : _GEN_240;
  assign _GEN_305 = 6'hf == _T_173 ? _GEN_4 : _GEN_241;
  assign _GEN_306 = 6'h10 == _T_173 ? _GEN_4 : _GEN_242;
  assign _GEN_307 = 6'h11 == _T_173 ? _GEN_4 : _GEN_243;
  assign _GEN_308 = 6'h12 == _T_173 ? _GEN_4 : _GEN_244;
  assign _GEN_309 = 6'h13 == _T_173 ? _GEN_4 : _GEN_245;
  assign _GEN_310 = 6'h14 == _T_173 ? _GEN_4 : _GEN_246;
  assign _GEN_311 = 6'h15 == _T_173 ? _GEN_4 : _GEN_247;
  assign _GEN_312 = 6'h16 == _T_173 ? _GEN_4 : _GEN_248;
  assign _GEN_313 = 6'h17 == _T_173 ? _GEN_4 : _GEN_249;
  assign _GEN_314 = 6'h18 == _T_173 ? _GEN_4 : _GEN_250;
  assign _GEN_315 = 6'h19 == _T_173 ? _GEN_4 : _GEN_251;
  assign _GEN_316 = 6'h1a == _T_173 ? _GEN_4 : _GEN_252;
  assign _GEN_317 = 6'h1b == _T_173 ? _GEN_4 : _GEN_253;
  assign _GEN_318 = 6'h1c == _T_173 ? _GEN_4 : _GEN_254;
  assign _GEN_319 = 6'h1d == _T_173 ? _GEN_4 : _GEN_255;
  assign _GEN_320 = 6'h1e == _T_173 ? _GEN_4 : _GEN_256;
  assign _GEN_321 = 6'h1f == _T_173 ? _GEN_4 : _GEN_257;
  assign _GEN_322 = 6'h20 == _T_173 ? _GEN_4 : _GEN_258;
  assign _GEN_323 = 6'h21 == _T_173 ? _GEN_4 : _GEN_259;
  assign _GEN_324 = 6'h22 == _T_173 ? _GEN_4 : _GEN_260;
  assign _GEN_325 = 6'h23 == _T_173 ? _GEN_4 : _GEN_261;
  assign _GEN_326 = 6'h24 == _T_173 ? _GEN_4 : _GEN_262;
  assign _GEN_327 = 6'h25 == _T_173 ? _GEN_4 : _GEN_263;
  assign _GEN_328 = 6'h26 == _T_173 ? _GEN_4 : _GEN_264;
  assign _GEN_329 = 6'h27 == _T_173 ? _GEN_4 : _GEN_265;
  assign _GEN_330 = 6'h28 == _T_173 ? _GEN_4 : _GEN_266;
  assign _GEN_331 = 6'h29 == _T_173 ? _GEN_4 : _GEN_267;
  assign _GEN_332 = 6'h2a == _T_173 ? _GEN_4 : _GEN_268;
  assign _GEN_333 = 6'h2b == _T_173 ? _GEN_4 : _GEN_269;
  assign _GEN_334 = 6'h2c == _T_173 ? _GEN_4 : _GEN_270;
  assign _GEN_335 = 6'h2d == _T_173 ? _GEN_4 : _GEN_271;
  assign _GEN_336 = 6'h2e == _T_173 ? _GEN_4 : _GEN_272;
  assign _GEN_337 = 6'h2f == _T_173 ? _GEN_4 : _GEN_273;
  assign _GEN_338 = 6'h30 == _T_173 ? _GEN_4 : _GEN_274;
  assign _GEN_339 = 6'h31 == _T_173 ? _GEN_4 : _GEN_275;
  assign _GEN_340 = 6'h32 == _T_173 ? _GEN_4 : _GEN_276;
  assign _GEN_341 = 6'h33 == _T_173 ? _GEN_4 : _GEN_277;
  assign _GEN_342 = 6'h34 == _T_173 ? _GEN_4 : _GEN_278;
  assign _GEN_343 = 6'h35 == _T_173 ? _GEN_4 : _GEN_279;
  assign _GEN_344 = 6'h36 == _T_173 ? _GEN_4 : _GEN_280;
  assign _GEN_345 = 6'h37 == _T_173 ? _GEN_4 : _GEN_281;
  assign _GEN_346 = 6'h38 == _T_173 ? _GEN_4 : _GEN_282;
  assign _GEN_347 = 6'h39 == _T_173 ? _GEN_4 : _GEN_283;
  assign _GEN_348 = 6'h3a == _T_173 ? _GEN_4 : _GEN_284;
  assign _GEN_349 = 6'h3b == _T_173 ? _GEN_4 : _GEN_285;
  assign _GEN_350 = 6'h3c == _T_173 ? _GEN_4 : _GEN_286;
  assign _GEN_351 = 6'h3d == _T_173 ? _GEN_4 : _GEN_287;
  assign _GEN_352 = 6'h3e == _T_173 ? _GEN_4 : _GEN_288;
  assign _GEN_353 = 6'h3f == _T_173 ? _GEN_4 : _GEN_289;
  assign _T_177 = wPos + 6'h5;
  assign _T_178 = _T_177[5:0];
  assign _T_180 = io_fastin[107:104];
  assign _GEN_5 = _T_180;
  assign _GEN_354 = 6'h0 == _T_178 ? _GEN_5 : _GEN_290;
  assign _GEN_355 = 6'h1 == _T_178 ? _GEN_5 : _GEN_291;
  assign _GEN_356 = 6'h2 == _T_178 ? _GEN_5 : _GEN_292;
  assign _GEN_357 = 6'h3 == _T_178 ? _GEN_5 : _GEN_293;
  assign _GEN_358 = 6'h4 == _T_178 ? _GEN_5 : _GEN_294;
  assign _GEN_359 = 6'h5 == _T_178 ? _GEN_5 : _GEN_295;
  assign _GEN_360 = 6'h6 == _T_178 ? _GEN_5 : _GEN_296;
  assign _GEN_361 = 6'h7 == _T_178 ? _GEN_5 : _GEN_297;
  assign _GEN_362 = 6'h8 == _T_178 ? _GEN_5 : _GEN_298;
  assign _GEN_363 = 6'h9 == _T_178 ? _GEN_5 : _GEN_299;
  assign _GEN_364 = 6'ha == _T_178 ? _GEN_5 : _GEN_300;
  assign _GEN_365 = 6'hb == _T_178 ? _GEN_5 : _GEN_301;
  assign _GEN_366 = 6'hc == _T_178 ? _GEN_5 : _GEN_302;
  assign _GEN_367 = 6'hd == _T_178 ? _GEN_5 : _GEN_303;
  assign _GEN_368 = 6'he == _T_178 ? _GEN_5 : _GEN_304;
  assign _GEN_369 = 6'hf == _T_178 ? _GEN_5 : _GEN_305;
  assign _GEN_370 = 6'h10 == _T_178 ? _GEN_5 : _GEN_306;
  assign _GEN_371 = 6'h11 == _T_178 ? _GEN_5 : _GEN_307;
  assign _GEN_372 = 6'h12 == _T_178 ? _GEN_5 : _GEN_308;
  assign _GEN_373 = 6'h13 == _T_178 ? _GEN_5 : _GEN_309;
  assign _GEN_374 = 6'h14 == _T_178 ? _GEN_5 : _GEN_310;
  assign _GEN_375 = 6'h15 == _T_178 ? _GEN_5 : _GEN_311;
  assign _GEN_376 = 6'h16 == _T_178 ? _GEN_5 : _GEN_312;
  assign _GEN_377 = 6'h17 == _T_178 ? _GEN_5 : _GEN_313;
  assign _GEN_378 = 6'h18 == _T_178 ? _GEN_5 : _GEN_314;
  assign _GEN_379 = 6'h19 == _T_178 ? _GEN_5 : _GEN_315;
  assign _GEN_380 = 6'h1a == _T_178 ? _GEN_5 : _GEN_316;
  assign _GEN_381 = 6'h1b == _T_178 ? _GEN_5 : _GEN_317;
  assign _GEN_382 = 6'h1c == _T_178 ? _GEN_5 : _GEN_318;
  assign _GEN_383 = 6'h1d == _T_178 ? _GEN_5 : _GEN_319;
  assign _GEN_384 = 6'h1e == _T_178 ? _GEN_5 : _GEN_320;
  assign _GEN_385 = 6'h1f == _T_178 ? _GEN_5 : _GEN_321;
  assign _GEN_386 = 6'h20 == _T_178 ? _GEN_5 : _GEN_322;
  assign _GEN_387 = 6'h21 == _T_178 ? _GEN_5 : _GEN_323;
  assign _GEN_388 = 6'h22 == _T_178 ? _GEN_5 : _GEN_324;
  assign _GEN_389 = 6'h23 == _T_178 ? _GEN_5 : _GEN_325;
  assign _GEN_390 = 6'h24 == _T_178 ? _GEN_5 : _GEN_326;
  assign _GEN_391 = 6'h25 == _T_178 ? _GEN_5 : _GEN_327;
  assign _GEN_392 = 6'h26 == _T_178 ? _GEN_5 : _GEN_328;
  assign _GEN_393 = 6'h27 == _T_178 ? _GEN_5 : _GEN_329;
  assign _GEN_394 = 6'h28 == _T_178 ? _GEN_5 : _GEN_330;
  assign _GEN_395 = 6'h29 == _T_178 ? _GEN_5 : _GEN_331;
  assign _GEN_396 = 6'h2a == _T_178 ? _GEN_5 : _GEN_332;
  assign _GEN_397 = 6'h2b == _T_178 ? _GEN_5 : _GEN_333;
  assign _GEN_398 = 6'h2c == _T_178 ? _GEN_5 : _GEN_334;
  assign _GEN_399 = 6'h2d == _T_178 ? _GEN_5 : _GEN_335;
  assign _GEN_400 = 6'h2e == _T_178 ? _GEN_5 : _GEN_336;
  assign _GEN_401 = 6'h2f == _T_178 ? _GEN_5 : _GEN_337;
  assign _GEN_402 = 6'h30 == _T_178 ? _GEN_5 : _GEN_338;
  assign _GEN_403 = 6'h31 == _T_178 ? _GEN_5 : _GEN_339;
  assign _GEN_404 = 6'h32 == _T_178 ? _GEN_5 : _GEN_340;
  assign _GEN_405 = 6'h33 == _T_178 ? _GEN_5 : _GEN_341;
  assign _GEN_406 = 6'h34 == _T_178 ? _GEN_5 : _GEN_342;
  assign _GEN_407 = 6'h35 == _T_178 ? _GEN_5 : _GEN_343;
  assign _GEN_408 = 6'h36 == _T_178 ? _GEN_5 : _GEN_344;
  assign _GEN_409 = 6'h37 == _T_178 ? _GEN_5 : _GEN_345;
  assign _GEN_410 = 6'h38 == _T_178 ? _GEN_5 : _GEN_346;
  assign _GEN_411 = 6'h39 == _T_178 ? _GEN_5 : _GEN_347;
  assign _GEN_412 = 6'h3a == _T_178 ? _GEN_5 : _GEN_348;
  assign _GEN_413 = 6'h3b == _T_178 ? _GEN_5 : _GEN_349;
  assign _GEN_414 = 6'h3c == _T_178 ? _GEN_5 : _GEN_350;
  assign _GEN_415 = 6'h3d == _T_178 ? _GEN_5 : _GEN_351;
  assign _GEN_416 = 6'h3e == _T_178 ? _GEN_5 : _GEN_352;
  assign _GEN_417 = 6'h3f == _T_178 ? _GEN_5 : _GEN_353;
  assign _T_182 = wPos + 6'h6;
  assign _T_183 = _T_182[5:0];
  assign _T_185 = io_fastin[103:100];
  assign _GEN_6 = _T_185;
  assign _GEN_418 = 6'h0 == _T_183 ? _GEN_6 : _GEN_354;
  assign _GEN_419 = 6'h1 == _T_183 ? _GEN_6 : _GEN_355;
  assign _GEN_420 = 6'h2 == _T_183 ? _GEN_6 : _GEN_356;
  assign _GEN_421 = 6'h3 == _T_183 ? _GEN_6 : _GEN_357;
  assign _GEN_422 = 6'h4 == _T_183 ? _GEN_6 : _GEN_358;
  assign _GEN_423 = 6'h5 == _T_183 ? _GEN_6 : _GEN_359;
  assign _GEN_424 = 6'h6 == _T_183 ? _GEN_6 : _GEN_360;
  assign _GEN_425 = 6'h7 == _T_183 ? _GEN_6 : _GEN_361;
  assign _GEN_426 = 6'h8 == _T_183 ? _GEN_6 : _GEN_362;
  assign _GEN_427 = 6'h9 == _T_183 ? _GEN_6 : _GEN_363;
  assign _GEN_428 = 6'ha == _T_183 ? _GEN_6 : _GEN_364;
  assign _GEN_429 = 6'hb == _T_183 ? _GEN_6 : _GEN_365;
  assign _GEN_430 = 6'hc == _T_183 ? _GEN_6 : _GEN_366;
  assign _GEN_431 = 6'hd == _T_183 ? _GEN_6 : _GEN_367;
  assign _GEN_432 = 6'he == _T_183 ? _GEN_6 : _GEN_368;
  assign _GEN_433 = 6'hf == _T_183 ? _GEN_6 : _GEN_369;
  assign _GEN_434 = 6'h10 == _T_183 ? _GEN_6 : _GEN_370;
  assign _GEN_435 = 6'h11 == _T_183 ? _GEN_6 : _GEN_371;
  assign _GEN_436 = 6'h12 == _T_183 ? _GEN_6 : _GEN_372;
  assign _GEN_437 = 6'h13 == _T_183 ? _GEN_6 : _GEN_373;
  assign _GEN_438 = 6'h14 == _T_183 ? _GEN_6 : _GEN_374;
  assign _GEN_439 = 6'h15 == _T_183 ? _GEN_6 : _GEN_375;
  assign _GEN_440 = 6'h16 == _T_183 ? _GEN_6 : _GEN_376;
  assign _GEN_441 = 6'h17 == _T_183 ? _GEN_6 : _GEN_377;
  assign _GEN_442 = 6'h18 == _T_183 ? _GEN_6 : _GEN_378;
  assign _GEN_443 = 6'h19 == _T_183 ? _GEN_6 : _GEN_379;
  assign _GEN_444 = 6'h1a == _T_183 ? _GEN_6 : _GEN_380;
  assign _GEN_445 = 6'h1b == _T_183 ? _GEN_6 : _GEN_381;
  assign _GEN_446 = 6'h1c == _T_183 ? _GEN_6 : _GEN_382;
  assign _GEN_447 = 6'h1d == _T_183 ? _GEN_6 : _GEN_383;
  assign _GEN_448 = 6'h1e == _T_183 ? _GEN_6 : _GEN_384;
  assign _GEN_449 = 6'h1f == _T_183 ? _GEN_6 : _GEN_385;
  assign _GEN_450 = 6'h20 == _T_183 ? _GEN_6 : _GEN_386;
  assign _GEN_451 = 6'h21 == _T_183 ? _GEN_6 : _GEN_387;
  assign _GEN_452 = 6'h22 == _T_183 ? _GEN_6 : _GEN_388;
  assign _GEN_453 = 6'h23 == _T_183 ? _GEN_6 : _GEN_389;
  assign _GEN_454 = 6'h24 == _T_183 ? _GEN_6 : _GEN_390;
  assign _GEN_455 = 6'h25 == _T_183 ? _GEN_6 : _GEN_391;
  assign _GEN_456 = 6'h26 == _T_183 ? _GEN_6 : _GEN_392;
  assign _GEN_457 = 6'h27 == _T_183 ? _GEN_6 : _GEN_393;
  assign _GEN_458 = 6'h28 == _T_183 ? _GEN_6 : _GEN_394;
  assign _GEN_459 = 6'h29 == _T_183 ? _GEN_6 : _GEN_395;
  assign _GEN_460 = 6'h2a == _T_183 ? _GEN_6 : _GEN_396;
  assign _GEN_461 = 6'h2b == _T_183 ? _GEN_6 : _GEN_397;
  assign _GEN_462 = 6'h2c == _T_183 ? _GEN_6 : _GEN_398;
  assign _GEN_463 = 6'h2d == _T_183 ? _GEN_6 : _GEN_399;
  assign _GEN_464 = 6'h2e == _T_183 ? _GEN_6 : _GEN_400;
  assign _GEN_465 = 6'h2f == _T_183 ? _GEN_6 : _GEN_401;
  assign _GEN_466 = 6'h30 == _T_183 ? _GEN_6 : _GEN_402;
  assign _GEN_467 = 6'h31 == _T_183 ? _GEN_6 : _GEN_403;
  assign _GEN_468 = 6'h32 == _T_183 ? _GEN_6 : _GEN_404;
  assign _GEN_469 = 6'h33 == _T_183 ? _GEN_6 : _GEN_405;
  assign _GEN_470 = 6'h34 == _T_183 ? _GEN_6 : _GEN_406;
  assign _GEN_471 = 6'h35 == _T_183 ? _GEN_6 : _GEN_407;
  assign _GEN_472 = 6'h36 == _T_183 ? _GEN_6 : _GEN_408;
  assign _GEN_473 = 6'h37 == _T_183 ? _GEN_6 : _GEN_409;
  assign _GEN_474 = 6'h38 == _T_183 ? _GEN_6 : _GEN_410;
  assign _GEN_475 = 6'h39 == _T_183 ? _GEN_6 : _GEN_411;
  assign _GEN_476 = 6'h3a == _T_183 ? _GEN_6 : _GEN_412;
  assign _GEN_477 = 6'h3b == _T_183 ? _GEN_6 : _GEN_413;
  assign _GEN_478 = 6'h3c == _T_183 ? _GEN_6 : _GEN_414;
  assign _GEN_479 = 6'h3d == _T_183 ? _GEN_6 : _GEN_415;
  assign _GEN_480 = 6'h3e == _T_183 ? _GEN_6 : _GEN_416;
  assign _GEN_481 = 6'h3f == _T_183 ? _GEN_6 : _GEN_417;
  assign _T_187 = wPos + 6'h7;
  assign _T_188 = _T_187[5:0];
  assign _T_190 = io_fastin[99:96];
  assign _GEN_7 = _T_190;
  assign _GEN_482 = 6'h0 == _T_188 ? _GEN_7 : _GEN_418;
  assign _GEN_483 = 6'h1 == _T_188 ? _GEN_7 : _GEN_419;
  assign _GEN_484 = 6'h2 == _T_188 ? _GEN_7 : _GEN_420;
  assign _GEN_485 = 6'h3 == _T_188 ? _GEN_7 : _GEN_421;
  assign _GEN_486 = 6'h4 == _T_188 ? _GEN_7 : _GEN_422;
  assign _GEN_487 = 6'h5 == _T_188 ? _GEN_7 : _GEN_423;
  assign _GEN_488 = 6'h6 == _T_188 ? _GEN_7 : _GEN_424;
  assign _GEN_489 = 6'h7 == _T_188 ? _GEN_7 : _GEN_425;
  assign _GEN_490 = 6'h8 == _T_188 ? _GEN_7 : _GEN_426;
  assign _GEN_491 = 6'h9 == _T_188 ? _GEN_7 : _GEN_427;
  assign _GEN_492 = 6'ha == _T_188 ? _GEN_7 : _GEN_428;
  assign _GEN_493 = 6'hb == _T_188 ? _GEN_7 : _GEN_429;
  assign _GEN_494 = 6'hc == _T_188 ? _GEN_7 : _GEN_430;
  assign _GEN_495 = 6'hd == _T_188 ? _GEN_7 : _GEN_431;
  assign _GEN_496 = 6'he == _T_188 ? _GEN_7 : _GEN_432;
  assign _GEN_497 = 6'hf == _T_188 ? _GEN_7 : _GEN_433;
  assign _GEN_498 = 6'h10 == _T_188 ? _GEN_7 : _GEN_434;
  assign _GEN_499 = 6'h11 == _T_188 ? _GEN_7 : _GEN_435;
  assign _GEN_500 = 6'h12 == _T_188 ? _GEN_7 : _GEN_436;
  assign _GEN_501 = 6'h13 == _T_188 ? _GEN_7 : _GEN_437;
  assign _GEN_502 = 6'h14 == _T_188 ? _GEN_7 : _GEN_438;
  assign _GEN_503 = 6'h15 == _T_188 ? _GEN_7 : _GEN_439;
  assign _GEN_504 = 6'h16 == _T_188 ? _GEN_7 : _GEN_440;
  assign _GEN_505 = 6'h17 == _T_188 ? _GEN_7 : _GEN_441;
  assign _GEN_506 = 6'h18 == _T_188 ? _GEN_7 : _GEN_442;
  assign _GEN_507 = 6'h19 == _T_188 ? _GEN_7 : _GEN_443;
  assign _GEN_508 = 6'h1a == _T_188 ? _GEN_7 : _GEN_444;
  assign _GEN_509 = 6'h1b == _T_188 ? _GEN_7 : _GEN_445;
  assign _GEN_510 = 6'h1c == _T_188 ? _GEN_7 : _GEN_446;
  assign _GEN_511 = 6'h1d == _T_188 ? _GEN_7 : _GEN_447;
  assign _GEN_512 = 6'h1e == _T_188 ? _GEN_7 : _GEN_448;
  assign _GEN_513 = 6'h1f == _T_188 ? _GEN_7 : _GEN_449;
  assign _GEN_514 = 6'h20 == _T_188 ? _GEN_7 : _GEN_450;
  assign _GEN_515 = 6'h21 == _T_188 ? _GEN_7 : _GEN_451;
  assign _GEN_516 = 6'h22 == _T_188 ? _GEN_7 : _GEN_452;
  assign _GEN_517 = 6'h23 == _T_188 ? _GEN_7 : _GEN_453;
  assign _GEN_518 = 6'h24 == _T_188 ? _GEN_7 : _GEN_454;
  assign _GEN_519 = 6'h25 == _T_188 ? _GEN_7 : _GEN_455;
  assign _GEN_520 = 6'h26 == _T_188 ? _GEN_7 : _GEN_456;
  assign _GEN_521 = 6'h27 == _T_188 ? _GEN_7 : _GEN_457;
  assign _GEN_522 = 6'h28 == _T_188 ? _GEN_7 : _GEN_458;
  assign _GEN_523 = 6'h29 == _T_188 ? _GEN_7 : _GEN_459;
  assign _GEN_524 = 6'h2a == _T_188 ? _GEN_7 : _GEN_460;
  assign _GEN_525 = 6'h2b == _T_188 ? _GEN_7 : _GEN_461;
  assign _GEN_526 = 6'h2c == _T_188 ? _GEN_7 : _GEN_462;
  assign _GEN_527 = 6'h2d == _T_188 ? _GEN_7 : _GEN_463;
  assign _GEN_528 = 6'h2e == _T_188 ? _GEN_7 : _GEN_464;
  assign _GEN_529 = 6'h2f == _T_188 ? _GEN_7 : _GEN_465;
  assign _GEN_530 = 6'h30 == _T_188 ? _GEN_7 : _GEN_466;
  assign _GEN_531 = 6'h31 == _T_188 ? _GEN_7 : _GEN_467;
  assign _GEN_532 = 6'h32 == _T_188 ? _GEN_7 : _GEN_468;
  assign _GEN_533 = 6'h33 == _T_188 ? _GEN_7 : _GEN_469;
  assign _GEN_534 = 6'h34 == _T_188 ? _GEN_7 : _GEN_470;
  assign _GEN_535 = 6'h35 == _T_188 ? _GEN_7 : _GEN_471;
  assign _GEN_536 = 6'h36 == _T_188 ? _GEN_7 : _GEN_472;
  assign _GEN_537 = 6'h37 == _T_188 ? _GEN_7 : _GEN_473;
  assign _GEN_538 = 6'h38 == _T_188 ? _GEN_7 : _GEN_474;
  assign _GEN_539 = 6'h39 == _T_188 ? _GEN_7 : _GEN_475;
  assign _GEN_540 = 6'h3a == _T_188 ? _GEN_7 : _GEN_476;
  assign _GEN_541 = 6'h3b == _T_188 ? _GEN_7 : _GEN_477;
  assign _GEN_542 = 6'h3c == _T_188 ? _GEN_7 : _GEN_478;
  assign _GEN_543 = 6'h3d == _T_188 ? _GEN_7 : _GEN_479;
  assign _GEN_544 = 6'h3e == _T_188 ? _GEN_7 : _GEN_480;
  assign _GEN_545 = 6'h3f == _T_188 ? _GEN_7 : _GEN_481;
  assign _T_192 = wPos + 6'h8;
  assign _T_193 = _T_192[5:0];
  assign _T_195 = io_fastin[95:92];
  assign _GEN_8 = _T_195;
  assign _GEN_546 = 6'h0 == _T_193 ? _GEN_8 : _GEN_482;
  assign _GEN_547 = 6'h1 == _T_193 ? _GEN_8 : _GEN_483;
  assign _GEN_548 = 6'h2 == _T_193 ? _GEN_8 : _GEN_484;
  assign _GEN_549 = 6'h3 == _T_193 ? _GEN_8 : _GEN_485;
  assign _GEN_550 = 6'h4 == _T_193 ? _GEN_8 : _GEN_486;
  assign _GEN_551 = 6'h5 == _T_193 ? _GEN_8 : _GEN_487;
  assign _GEN_552 = 6'h6 == _T_193 ? _GEN_8 : _GEN_488;
  assign _GEN_553 = 6'h7 == _T_193 ? _GEN_8 : _GEN_489;
  assign _GEN_554 = 6'h8 == _T_193 ? _GEN_8 : _GEN_490;
  assign _GEN_555 = 6'h9 == _T_193 ? _GEN_8 : _GEN_491;
  assign _GEN_556 = 6'ha == _T_193 ? _GEN_8 : _GEN_492;
  assign _GEN_557 = 6'hb == _T_193 ? _GEN_8 : _GEN_493;
  assign _GEN_558 = 6'hc == _T_193 ? _GEN_8 : _GEN_494;
  assign _GEN_559 = 6'hd == _T_193 ? _GEN_8 : _GEN_495;
  assign _GEN_560 = 6'he == _T_193 ? _GEN_8 : _GEN_496;
  assign _GEN_561 = 6'hf == _T_193 ? _GEN_8 : _GEN_497;
  assign _GEN_562 = 6'h10 == _T_193 ? _GEN_8 : _GEN_498;
  assign _GEN_563 = 6'h11 == _T_193 ? _GEN_8 : _GEN_499;
  assign _GEN_564 = 6'h12 == _T_193 ? _GEN_8 : _GEN_500;
  assign _GEN_565 = 6'h13 == _T_193 ? _GEN_8 : _GEN_501;
  assign _GEN_566 = 6'h14 == _T_193 ? _GEN_8 : _GEN_502;
  assign _GEN_567 = 6'h15 == _T_193 ? _GEN_8 : _GEN_503;
  assign _GEN_568 = 6'h16 == _T_193 ? _GEN_8 : _GEN_504;
  assign _GEN_569 = 6'h17 == _T_193 ? _GEN_8 : _GEN_505;
  assign _GEN_570 = 6'h18 == _T_193 ? _GEN_8 : _GEN_506;
  assign _GEN_571 = 6'h19 == _T_193 ? _GEN_8 : _GEN_507;
  assign _GEN_572 = 6'h1a == _T_193 ? _GEN_8 : _GEN_508;
  assign _GEN_573 = 6'h1b == _T_193 ? _GEN_8 : _GEN_509;
  assign _GEN_574 = 6'h1c == _T_193 ? _GEN_8 : _GEN_510;
  assign _GEN_575 = 6'h1d == _T_193 ? _GEN_8 : _GEN_511;
  assign _GEN_576 = 6'h1e == _T_193 ? _GEN_8 : _GEN_512;
  assign _GEN_577 = 6'h1f == _T_193 ? _GEN_8 : _GEN_513;
  assign _GEN_578 = 6'h20 == _T_193 ? _GEN_8 : _GEN_514;
  assign _GEN_579 = 6'h21 == _T_193 ? _GEN_8 : _GEN_515;
  assign _GEN_580 = 6'h22 == _T_193 ? _GEN_8 : _GEN_516;
  assign _GEN_581 = 6'h23 == _T_193 ? _GEN_8 : _GEN_517;
  assign _GEN_582 = 6'h24 == _T_193 ? _GEN_8 : _GEN_518;
  assign _GEN_583 = 6'h25 == _T_193 ? _GEN_8 : _GEN_519;
  assign _GEN_584 = 6'h26 == _T_193 ? _GEN_8 : _GEN_520;
  assign _GEN_585 = 6'h27 == _T_193 ? _GEN_8 : _GEN_521;
  assign _GEN_586 = 6'h28 == _T_193 ? _GEN_8 : _GEN_522;
  assign _GEN_587 = 6'h29 == _T_193 ? _GEN_8 : _GEN_523;
  assign _GEN_588 = 6'h2a == _T_193 ? _GEN_8 : _GEN_524;
  assign _GEN_589 = 6'h2b == _T_193 ? _GEN_8 : _GEN_525;
  assign _GEN_590 = 6'h2c == _T_193 ? _GEN_8 : _GEN_526;
  assign _GEN_591 = 6'h2d == _T_193 ? _GEN_8 : _GEN_527;
  assign _GEN_592 = 6'h2e == _T_193 ? _GEN_8 : _GEN_528;
  assign _GEN_593 = 6'h2f == _T_193 ? _GEN_8 : _GEN_529;
  assign _GEN_594 = 6'h30 == _T_193 ? _GEN_8 : _GEN_530;
  assign _GEN_595 = 6'h31 == _T_193 ? _GEN_8 : _GEN_531;
  assign _GEN_596 = 6'h32 == _T_193 ? _GEN_8 : _GEN_532;
  assign _GEN_597 = 6'h33 == _T_193 ? _GEN_8 : _GEN_533;
  assign _GEN_598 = 6'h34 == _T_193 ? _GEN_8 : _GEN_534;
  assign _GEN_599 = 6'h35 == _T_193 ? _GEN_8 : _GEN_535;
  assign _GEN_600 = 6'h36 == _T_193 ? _GEN_8 : _GEN_536;
  assign _GEN_601 = 6'h37 == _T_193 ? _GEN_8 : _GEN_537;
  assign _GEN_602 = 6'h38 == _T_193 ? _GEN_8 : _GEN_538;
  assign _GEN_603 = 6'h39 == _T_193 ? _GEN_8 : _GEN_539;
  assign _GEN_604 = 6'h3a == _T_193 ? _GEN_8 : _GEN_540;
  assign _GEN_605 = 6'h3b == _T_193 ? _GEN_8 : _GEN_541;
  assign _GEN_606 = 6'h3c == _T_193 ? _GEN_8 : _GEN_542;
  assign _GEN_607 = 6'h3d == _T_193 ? _GEN_8 : _GEN_543;
  assign _GEN_608 = 6'h3e == _T_193 ? _GEN_8 : _GEN_544;
  assign _GEN_609 = 6'h3f == _T_193 ? _GEN_8 : _GEN_545;
  assign _T_197 = wPos + 6'h9;
  assign _T_198 = _T_197[5:0];
  assign _T_200 = io_fastin[91:88];
  assign _GEN_9 = _T_200;
  assign _GEN_610 = 6'h0 == _T_198 ? _GEN_9 : _GEN_546;
  assign _GEN_611 = 6'h1 == _T_198 ? _GEN_9 : _GEN_547;
  assign _GEN_612 = 6'h2 == _T_198 ? _GEN_9 : _GEN_548;
  assign _GEN_613 = 6'h3 == _T_198 ? _GEN_9 : _GEN_549;
  assign _GEN_614 = 6'h4 == _T_198 ? _GEN_9 : _GEN_550;
  assign _GEN_615 = 6'h5 == _T_198 ? _GEN_9 : _GEN_551;
  assign _GEN_616 = 6'h6 == _T_198 ? _GEN_9 : _GEN_552;
  assign _GEN_617 = 6'h7 == _T_198 ? _GEN_9 : _GEN_553;
  assign _GEN_618 = 6'h8 == _T_198 ? _GEN_9 : _GEN_554;
  assign _GEN_619 = 6'h9 == _T_198 ? _GEN_9 : _GEN_555;
  assign _GEN_620 = 6'ha == _T_198 ? _GEN_9 : _GEN_556;
  assign _GEN_621 = 6'hb == _T_198 ? _GEN_9 : _GEN_557;
  assign _GEN_622 = 6'hc == _T_198 ? _GEN_9 : _GEN_558;
  assign _GEN_623 = 6'hd == _T_198 ? _GEN_9 : _GEN_559;
  assign _GEN_624 = 6'he == _T_198 ? _GEN_9 : _GEN_560;
  assign _GEN_625 = 6'hf == _T_198 ? _GEN_9 : _GEN_561;
  assign _GEN_626 = 6'h10 == _T_198 ? _GEN_9 : _GEN_562;
  assign _GEN_627 = 6'h11 == _T_198 ? _GEN_9 : _GEN_563;
  assign _GEN_628 = 6'h12 == _T_198 ? _GEN_9 : _GEN_564;
  assign _GEN_629 = 6'h13 == _T_198 ? _GEN_9 : _GEN_565;
  assign _GEN_630 = 6'h14 == _T_198 ? _GEN_9 : _GEN_566;
  assign _GEN_631 = 6'h15 == _T_198 ? _GEN_9 : _GEN_567;
  assign _GEN_632 = 6'h16 == _T_198 ? _GEN_9 : _GEN_568;
  assign _GEN_633 = 6'h17 == _T_198 ? _GEN_9 : _GEN_569;
  assign _GEN_634 = 6'h18 == _T_198 ? _GEN_9 : _GEN_570;
  assign _GEN_635 = 6'h19 == _T_198 ? _GEN_9 : _GEN_571;
  assign _GEN_636 = 6'h1a == _T_198 ? _GEN_9 : _GEN_572;
  assign _GEN_637 = 6'h1b == _T_198 ? _GEN_9 : _GEN_573;
  assign _GEN_638 = 6'h1c == _T_198 ? _GEN_9 : _GEN_574;
  assign _GEN_639 = 6'h1d == _T_198 ? _GEN_9 : _GEN_575;
  assign _GEN_640 = 6'h1e == _T_198 ? _GEN_9 : _GEN_576;
  assign _GEN_641 = 6'h1f == _T_198 ? _GEN_9 : _GEN_577;
  assign _GEN_642 = 6'h20 == _T_198 ? _GEN_9 : _GEN_578;
  assign _GEN_643 = 6'h21 == _T_198 ? _GEN_9 : _GEN_579;
  assign _GEN_644 = 6'h22 == _T_198 ? _GEN_9 : _GEN_580;
  assign _GEN_645 = 6'h23 == _T_198 ? _GEN_9 : _GEN_581;
  assign _GEN_646 = 6'h24 == _T_198 ? _GEN_9 : _GEN_582;
  assign _GEN_647 = 6'h25 == _T_198 ? _GEN_9 : _GEN_583;
  assign _GEN_648 = 6'h26 == _T_198 ? _GEN_9 : _GEN_584;
  assign _GEN_649 = 6'h27 == _T_198 ? _GEN_9 : _GEN_585;
  assign _GEN_650 = 6'h28 == _T_198 ? _GEN_9 : _GEN_586;
  assign _GEN_651 = 6'h29 == _T_198 ? _GEN_9 : _GEN_587;
  assign _GEN_652 = 6'h2a == _T_198 ? _GEN_9 : _GEN_588;
  assign _GEN_653 = 6'h2b == _T_198 ? _GEN_9 : _GEN_589;
  assign _GEN_654 = 6'h2c == _T_198 ? _GEN_9 : _GEN_590;
  assign _GEN_655 = 6'h2d == _T_198 ? _GEN_9 : _GEN_591;
  assign _GEN_656 = 6'h2e == _T_198 ? _GEN_9 : _GEN_592;
  assign _GEN_657 = 6'h2f == _T_198 ? _GEN_9 : _GEN_593;
  assign _GEN_658 = 6'h30 == _T_198 ? _GEN_9 : _GEN_594;
  assign _GEN_659 = 6'h31 == _T_198 ? _GEN_9 : _GEN_595;
  assign _GEN_660 = 6'h32 == _T_198 ? _GEN_9 : _GEN_596;
  assign _GEN_661 = 6'h33 == _T_198 ? _GEN_9 : _GEN_597;
  assign _GEN_662 = 6'h34 == _T_198 ? _GEN_9 : _GEN_598;
  assign _GEN_663 = 6'h35 == _T_198 ? _GEN_9 : _GEN_599;
  assign _GEN_664 = 6'h36 == _T_198 ? _GEN_9 : _GEN_600;
  assign _GEN_665 = 6'h37 == _T_198 ? _GEN_9 : _GEN_601;
  assign _GEN_666 = 6'h38 == _T_198 ? _GEN_9 : _GEN_602;
  assign _GEN_667 = 6'h39 == _T_198 ? _GEN_9 : _GEN_603;
  assign _GEN_668 = 6'h3a == _T_198 ? _GEN_9 : _GEN_604;
  assign _GEN_669 = 6'h3b == _T_198 ? _GEN_9 : _GEN_605;
  assign _GEN_670 = 6'h3c == _T_198 ? _GEN_9 : _GEN_606;
  assign _GEN_671 = 6'h3d == _T_198 ? _GEN_9 : _GEN_607;
  assign _GEN_672 = 6'h3e == _T_198 ? _GEN_9 : _GEN_608;
  assign _GEN_673 = 6'h3f == _T_198 ? _GEN_9 : _GEN_609;
  assign _T_202 = wPos + 6'ha;
  assign _T_203 = _T_202[5:0];
  assign _T_205 = io_fastin[87:84];
  assign _GEN_10 = _T_205;
  assign _GEN_674 = 6'h0 == _T_203 ? _GEN_10 : _GEN_610;
  assign _GEN_675 = 6'h1 == _T_203 ? _GEN_10 : _GEN_611;
  assign _GEN_676 = 6'h2 == _T_203 ? _GEN_10 : _GEN_612;
  assign _GEN_677 = 6'h3 == _T_203 ? _GEN_10 : _GEN_613;
  assign _GEN_678 = 6'h4 == _T_203 ? _GEN_10 : _GEN_614;
  assign _GEN_679 = 6'h5 == _T_203 ? _GEN_10 : _GEN_615;
  assign _GEN_680 = 6'h6 == _T_203 ? _GEN_10 : _GEN_616;
  assign _GEN_681 = 6'h7 == _T_203 ? _GEN_10 : _GEN_617;
  assign _GEN_682 = 6'h8 == _T_203 ? _GEN_10 : _GEN_618;
  assign _GEN_683 = 6'h9 == _T_203 ? _GEN_10 : _GEN_619;
  assign _GEN_684 = 6'ha == _T_203 ? _GEN_10 : _GEN_620;
  assign _GEN_685 = 6'hb == _T_203 ? _GEN_10 : _GEN_621;
  assign _GEN_686 = 6'hc == _T_203 ? _GEN_10 : _GEN_622;
  assign _GEN_687 = 6'hd == _T_203 ? _GEN_10 : _GEN_623;
  assign _GEN_688 = 6'he == _T_203 ? _GEN_10 : _GEN_624;
  assign _GEN_689 = 6'hf == _T_203 ? _GEN_10 : _GEN_625;
  assign _GEN_690 = 6'h10 == _T_203 ? _GEN_10 : _GEN_626;
  assign _GEN_691 = 6'h11 == _T_203 ? _GEN_10 : _GEN_627;
  assign _GEN_692 = 6'h12 == _T_203 ? _GEN_10 : _GEN_628;
  assign _GEN_693 = 6'h13 == _T_203 ? _GEN_10 : _GEN_629;
  assign _GEN_694 = 6'h14 == _T_203 ? _GEN_10 : _GEN_630;
  assign _GEN_695 = 6'h15 == _T_203 ? _GEN_10 : _GEN_631;
  assign _GEN_696 = 6'h16 == _T_203 ? _GEN_10 : _GEN_632;
  assign _GEN_697 = 6'h17 == _T_203 ? _GEN_10 : _GEN_633;
  assign _GEN_698 = 6'h18 == _T_203 ? _GEN_10 : _GEN_634;
  assign _GEN_699 = 6'h19 == _T_203 ? _GEN_10 : _GEN_635;
  assign _GEN_700 = 6'h1a == _T_203 ? _GEN_10 : _GEN_636;
  assign _GEN_701 = 6'h1b == _T_203 ? _GEN_10 : _GEN_637;
  assign _GEN_702 = 6'h1c == _T_203 ? _GEN_10 : _GEN_638;
  assign _GEN_703 = 6'h1d == _T_203 ? _GEN_10 : _GEN_639;
  assign _GEN_704 = 6'h1e == _T_203 ? _GEN_10 : _GEN_640;
  assign _GEN_705 = 6'h1f == _T_203 ? _GEN_10 : _GEN_641;
  assign _GEN_706 = 6'h20 == _T_203 ? _GEN_10 : _GEN_642;
  assign _GEN_707 = 6'h21 == _T_203 ? _GEN_10 : _GEN_643;
  assign _GEN_708 = 6'h22 == _T_203 ? _GEN_10 : _GEN_644;
  assign _GEN_709 = 6'h23 == _T_203 ? _GEN_10 : _GEN_645;
  assign _GEN_710 = 6'h24 == _T_203 ? _GEN_10 : _GEN_646;
  assign _GEN_711 = 6'h25 == _T_203 ? _GEN_10 : _GEN_647;
  assign _GEN_712 = 6'h26 == _T_203 ? _GEN_10 : _GEN_648;
  assign _GEN_713 = 6'h27 == _T_203 ? _GEN_10 : _GEN_649;
  assign _GEN_714 = 6'h28 == _T_203 ? _GEN_10 : _GEN_650;
  assign _GEN_715 = 6'h29 == _T_203 ? _GEN_10 : _GEN_651;
  assign _GEN_716 = 6'h2a == _T_203 ? _GEN_10 : _GEN_652;
  assign _GEN_717 = 6'h2b == _T_203 ? _GEN_10 : _GEN_653;
  assign _GEN_718 = 6'h2c == _T_203 ? _GEN_10 : _GEN_654;
  assign _GEN_719 = 6'h2d == _T_203 ? _GEN_10 : _GEN_655;
  assign _GEN_720 = 6'h2e == _T_203 ? _GEN_10 : _GEN_656;
  assign _GEN_721 = 6'h2f == _T_203 ? _GEN_10 : _GEN_657;
  assign _GEN_722 = 6'h30 == _T_203 ? _GEN_10 : _GEN_658;
  assign _GEN_723 = 6'h31 == _T_203 ? _GEN_10 : _GEN_659;
  assign _GEN_724 = 6'h32 == _T_203 ? _GEN_10 : _GEN_660;
  assign _GEN_725 = 6'h33 == _T_203 ? _GEN_10 : _GEN_661;
  assign _GEN_726 = 6'h34 == _T_203 ? _GEN_10 : _GEN_662;
  assign _GEN_727 = 6'h35 == _T_203 ? _GEN_10 : _GEN_663;
  assign _GEN_728 = 6'h36 == _T_203 ? _GEN_10 : _GEN_664;
  assign _GEN_729 = 6'h37 == _T_203 ? _GEN_10 : _GEN_665;
  assign _GEN_730 = 6'h38 == _T_203 ? _GEN_10 : _GEN_666;
  assign _GEN_731 = 6'h39 == _T_203 ? _GEN_10 : _GEN_667;
  assign _GEN_732 = 6'h3a == _T_203 ? _GEN_10 : _GEN_668;
  assign _GEN_733 = 6'h3b == _T_203 ? _GEN_10 : _GEN_669;
  assign _GEN_734 = 6'h3c == _T_203 ? _GEN_10 : _GEN_670;
  assign _GEN_735 = 6'h3d == _T_203 ? _GEN_10 : _GEN_671;
  assign _GEN_736 = 6'h3e == _T_203 ? _GEN_10 : _GEN_672;
  assign _GEN_737 = 6'h3f == _T_203 ? _GEN_10 : _GEN_673;
  assign _T_207 = wPos + 6'hb;
  assign _T_208 = _T_207[5:0];
  assign _T_210 = io_fastin[83:80];
  assign _GEN_11 = _T_210;
  assign _GEN_738 = 6'h0 == _T_208 ? _GEN_11 : _GEN_674;
  assign _GEN_739 = 6'h1 == _T_208 ? _GEN_11 : _GEN_675;
  assign _GEN_740 = 6'h2 == _T_208 ? _GEN_11 : _GEN_676;
  assign _GEN_741 = 6'h3 == _T_208 ? _GEN_11 : _GEN_677;
  assign _GEN_742 = 6'h4 == _T_208 ? _GEN_11 : _GEN_678;
  assign _GEN_743 = 6'h5 == _T_208 ? _GEN_11 : _GEN_679;
  assign _GEN_744 = 6'h6 == _T_208 ? _GEN_11 : _GEN_680;
  assign _GEN_745 = 6'h7 == _T_208 ? _GEN_11 : _GEN_681;
  assign _GEN_746 = 6'h8 == _T_208 ? _GEN_11 : _GEN_682;
  assign _GEN_747 = 6'h9 == _T_208 ? _GEN_11 : _GEN_683;
  assign _GEN_748 = 6'ha == _T_208 ? _GEN_11 : _GEN_684;
  assign _GEN_749 = 6'hb == _T_208 ? _GEN_11 : _GEN_685;
  assign _GEN_750 = 6'hc == _T_208 ? _GEN_11 : _GEN_686;
  assign _GEN_751 = 6'hd == _T_208 ? _GEN_11 : _GEN_687;
  assign _GEN_752 = 6'he == _T_208 ? _GEN_11 : _GEN_688;
  assign _GEN_753 = 6'hf == _T_208 ? _GEN_11 : _GEN_689;
  assign _GEN_754 = 6'h10 == _T_208 ? _GEN_11 : _GEN_690;
  assign _GEN_755 = 6'h11 == _T_208 ? _GEN_11 : _GEN_691;
  assign _GEN_756 = 6'h12 == _T_208 ? _GEN_11 : _GEN_692;
  assign _GEN_757 = 6'h13 == _T_208 ? _GEN_11 : _GEN_693;
  assign _GEN_758 = 6'h14 == _T_208 ? _GEN_11 : _GEN_694;
  assign _GEN_759 = 6'h15 == _T_208 ? _GEN_11 : _GEN_695;
  assign _GEN_760 = 6'h16 == _T_208 ? _GEN_11 : _GEN_696;
  assign _GEN_761 = 6'h17 == _T_208 ? _GEN_11 : _GEN_697;
  assign _GEN_762 = 6'h18 == _T_208 ? _GEN_11 : _GEN_698;
  assign _GEN_763 = 6'h19 == _T_208 ? _GEN_11 : _GEN_699;
  assign _GEN_764 = 6'h1a == _T_208 ? _GEN_11 : _GEN_700;
  assign _GEN_765 = 6'h1b == _T_208 ? _GEN_11 : _GEN_701;
  assign _GEN_766 = 6'h1c == _T_208 ? _GEN_11 : _GEN_702;
  assign _GEN_767 = 6'h1d == _T_208 ? _GEN_11 : _GEN_703;
  assign _GEN_768 = 6'h1e == _T_208 ? _GEN_11 : _GEN_704;
  assign _GEN_769 = 6'h1f == _T_208 ? _GEN_11 : _GEN_705;
  assign _GEN_770 = 6'h20 == _T_208 ? _GEN_11 : _GEN_706;
  assign _GEN_771 = 6'h21 == _T_208 ? _GEN_11 : _GEN_707;
  assign _GEN_772 = 6'h22 == _T_208 ? _GEN_11 : _GEN_708;
  assign _GEN_773 = 6'h23 == _T_208 ? _GEN_11 : _GEN_709;
  assign _GEN_774 = 6'h24 == _T_208 ? _GEN_11 : _GEN_710;
  assign _GEN_775 = 6'h25 == _T_208 ? _GEN_11 : _GEN_711;
  assign _GEN_776 = 6'h26 == _T_208 ? _GEN_11 : _GEN_712;
  assign _GEN_777 = 6'h27 == _T_208 ? _GEN_11 : _GEN_713;
  assign _GEN_778 = 6'h28 == _T_208 ? _GEN_11 : _GEN_714;
  assign _GEN_779 = 6'h29 == _T_208 ? _GEN_11 : _GEN_715;
  assign _GEN_780 = 6'h2a == _T_208 ? _GEN_11 : _GEN_716;
  assign _GEN_781 = 6'h2b == _T_208 ? _GEN_11 : _GEN_717;
  assign _GEN_782 = 6'h2c == _T_208 ? _GEN_11 : _GEN_718;
  assign _GEN_783 = 6'h2d == _T_208 ? _GEN_11 : _GEN_719;
  assign _GEN_784 = 6'h2e == _T_208 ? _GEN_11 : _GEN_720;
  assign _GEN_785 = 6'h2f == _T_208 ? _GEN_11 : _GEN_721;
  assign _GEN_786 = 6'h30 == _T_208 ? _GEN_11 : _GEN_722;
  assign _GEN_787 = 6'h31 == _T_208 ? _GEN_11 : _GEN_723;
  assign _GEN_788 = 6'h32 == _T_208 ? _GEN_11 : _GEN_724;
  assign _GEN_789 = 6'h33 == _T_208 ? _GEN_11 : _GEN_725;
  assign _GEN_790 = 6'h34 == _T_208 ? _GEN_11 : _GEN_726;
  assign _GEN_791 = 6'h35 == _T_208 ? _GEN_11 : _GEN_727;
  assign _GEN_792 = 6'h36 == _T_208 ? _GEN_11 : _GEN_728;
  assign _GEN_793 = 6'h37 == _T_208 ? _GEN_11 : _GEN_729;
  assign _GEN_794 = 6'h38 == _T_208 ? _GEN_11 : _GEN_730;
  assign _GEN_795 = 6'h39 == _T_208 ? _GEN_11 : _GEN_731;
  assign _GEN_796 = 6'h3a == _T_208 ? _GEN_11 : _GEN_732;
  assign _GEN_797 = 6'h3b == _T_208 ? _GEN_11 : _GEN_733;
  assign _GEN_798 = 6'h3c == _T_208 ? _GEN_11 : _GEN_734;
  assign _GEN_799 = 6'h3d == _T_208 ? _GEN_11 : _GEN_735;
  assign _GEN_800 = 6'h3e == _T_208 ? _GEN_11 : _GEN_736;
  assign _GEN_801 = 6'h3f == _T_208 ? _GEN_11 : _GEN_737;
  assign _T_212 = wPos + 6'hc;
  assign _T_213 = _T_212[5:0];
  assign _T_215 = io_fastin[79:76];
  assign _GEN_12 = _T_215;
  assign _GEN_802 = 6'h0 == _T_213 ? _GEN_12 : _GEN_738;
  assign _GEN_803 = 6'h1 == _T_213 ? _GEN_12 : _GEN_739;
  assign _GEN_804 = 6'h2 == _T_213 ? _GEN_12 : _GEN_740;
  assign _GEN_805 = 6'h3 == _T_213 ? _GEN_12 : _GEN_741;
  assign _GEN_806 = 6'h4 == _T_213 ? _GEN_12 : _GEN_742;
  assign _GEN_807 = 6'h5 == _T_213 ? _GEN_12 : _GEN_743;
  assign _GEN_808 = 6'h6 == _T_213 ? _GEN_12 : _GEN_744;
  assign _GEN_809 = 6'h7 == _T_213 ? _GEN_12 : _GEN_745;
  assign _GEN_810 = 6'h8 == _T_213 ? _GEN_12 : _GEN_746;
  assign _GEN_811 = 6'h9 == _T_213 ? _GEN_12 : _GEN_747;
  assign _GEN_812 = 6'ha == _T_213 ? _GEN_12 : _GEN_748;
  assign _GEN_813 = 6'hb == _T_213 ? _GEN_12 : _GEN_749;
  assign _GEN_814 = 6'hc == _T_213 ? _GEN_12 : _GEN_750;
  assign _GEN_815 = 6'hd == _T_213 ? _GEN_12 : _GEN_751;
  assign _GEN_816 = 6'he == _T_213 ? _GEN_12 : _GEN_752;
  assign _GEN_817 = 6'hf == _T_213 ? _GEN_12 : _GEN_753;
  assign _GEN_818 = 6'h10 == _T_213 ? _GEN_12 : _GEN_754;
  assign _GEN_819 = 6'h11 == _T_213 ? _GEN_12 : _GEN_755;
  assign _GEN_820 = 6'h12 == _T_213 ? _GEN_12 : _GEN_756;
  assign _GEN_821 = 6'h13 == _T_213 ? _GEN_12 : _GEN_757;
  assign _GEN_822 = 6'h14 == _T_213 ? _GEN_12 : _GEN_758;
  assign _GEN_823 = 6'h15 == _T_213 ? _GEN_12 : _GEN_759;
  assign _GEN_824 = 6'h16 == _T_213 ? _GEN_12 : _GEN_760;
  assign _GEN_825 = 6'h17 == _T_213 ? _GEN_12 : _GEN_761;
  assign _GEN_826 = 6'h18 == _T_213 ? _GEN_12 : _GEN_762;
  assign _GEN_827 = 6'h19 == _T_213 ? _GEN_12 : _GEN_763;
  assign _GEN_828 = 6'h1a == _T_213 ? _GEN_12 : _GEN_764;
  assign _GEN_829 = 6'h1b == _T_213 ? _GEN_12 : _GEN_765;
  assign _GEN_830 = 6'h1c == _T_213 ? _GEN_12 : _GEN_766;
  assign _GEN_831 = 6'h1d == _T_213 ? _GEN_12 : _GEN_767;
  assign _GEN_832 = 6'h1e == _T_213 ? _GEN_12 : _GEN_768;
  assign _GEN_833 = 6'h1f == _T_213 ? _GEN_12 : _GEN_769;
  assign _GEN_834 = 6'h20 == _T_213 ? _GEN_12 : _GEN_770;
  assign _GEN_835 = 6'h21 == _T_213 ? _GEN_12 : _GEN_771;
  assign _GEN_836 = 6'h22 == _T_213 ? _GEN_12 : _GEN_772;
  assign _GEN_837 = 6'h23 == _T_213 ? _GEN_12 : _GEN_773;
  assign _GEN_838 = 6'h24 == _T_213 ? _GEN_12 : _GEN_774;
  assign _GEN_839 = 6'h25 == _T_213 ? _GEN_12 : _GEN_775;
  assign _GEN_840 = 6'h26 == _T_213 ? _GEN_12 : _GEN_776;
  assign _GEN_841 = 6'h27 == _T_213 ? _GEN_12 : _GEN_777;
  assign _GEN_842 = 6'h28 == _T_213 ? _GEN_12 : _GEN_778;
  assign _GEN_843 = 6'h29 == _T_213 ? _GEN_12 : _GEN_779;
  assign _GEN_844 = 6'h2a == _T_213 ? _GEN_12 : _GEN_780;
  assign _GEN_845 = 6'h2b == _T_213 ? _GEN_12 : _GEN_781;
  assign _GEN_846 = 6'h2c == _T_213 ? _GEN_12 : _GEN_782;
  assign _GEN_847 = 6'h2d == _T_213 ? _GEN_12 : _GEN_783;
  assign _GEN_848 = 6'h2e == _T_213 ? _GEN_12 : _GEN_784;
  assign _GEN_849 = 6'h2f == _T_213 ? _GEN_12 : _GEN_785;
  assign _GEN_850 = 6'h30 == _T_213 ? _GEN_12 : _GEN_786;
  assign _GEN_851 = 6'h31 == _T_213 ? _GEN_12 : _GEN_787;
  assign _GEN_852 = 6'h32 == _T_213 ? _GEN_12 : _GEN_788;
  assign _GEN_853 = 6'h33 == _T_213 ? _GEN_12 : _GEN_789;
  assign _GEN_854 = 6'h34 == _T_213 ? _GEN_12 : _GEN_790;
  assign _GEN_855 = 6'h35 == _T_213 ? _GEN_12 : _GEN_791;
  assign _GEN_856 = 6'h36 == _T_213 ? _GEN_12 : _GEN_792;
  assign _GEN_857 = 6'h37 == _T_213 ? _GEN_12 : _GEN_793;
  assign _GEN_858 = 6'h38 == _T_213 ? _GEN_12 : _GEN_794;
  assign _GEN_859 = 6'h39 == _T_213 ? _GEN_12 : _GEN_795;
  assign _GEN_860 = 6'h3a == _T_213 ? _GEN_12 : _GEN_796;
  assign _GEN_861 = 6'h3b == _T_213 ? _GEN_12 : _GEN_797;
  assign _GEN_862 = 6'h3c == _T_213 ? _GEN_12 : _GEN_798;
  assign _GEN_863 = 6'h3d == _T_213 ? _GEN_12 : _GEN_799;
  assign _GEN_864 = 6'h3e == _T_213 ? _GEN_12 : _GEN_800;
  assign _GEN_865 = 6'h3f == _T_213 ? _GEN_12 : _GEN_801;
  assign _T_217 = wPos + 6'hd;
  assign _T_218 = _T_217[5:0];
  assign _T_220 = io_fastin[75:72];
  assign _GEN_13 = _T_220;
  assign _GEN_866 = 6'h0 == _T_218 ? _GEN_13 : _GEN_802;
  assign _GEN_867 = 6'h1 == _T_218 ? _GEN_13 : _GEN_803;
  assign _GEN_868 = 6'h2 == _T_218 ? _GEN_13 : _GEN_804;
  assign _GEN_869 = 6'h3 == _T_218 ? _GEN_13 : _GEN_805;
  assign _GEN_870 = 6'h4 == _T_218 ? _GEN_13 : _GEN_806;
  assign _GEN_871 = 6'h5 == _T_218 ? _GEN_13 : _GEN_807;
  assign _GEN_872 = 6'h6 == _T_218 ? _GEN_13 : _GEN_808;
  assign _GEN_873 = 6'h7 == _T_218 ? _GEN_13 : _GEN_809;
  assign _GEN_874 = 6'h8 == _T_218 ? _GEN_13 : _GEN_810;
  assign _GEN_875 = 6'h9 == _T_218 ? _GEN_13 : _GEN_811;
  assign _GEN_876 = 6'ha == _T_218 ? _GEN_13 : _GEN_812;
  assign _GEN_877 = 6'hb == _T_218 ? _GEN_13 : _GEN_813;
  assign _GEN_878 = 6'hc == _T_218 ? _GEN_13 : _GEN_814;
  assign _GEN_879 = 6'hd == _T_218 ? _GEN_13 : _GEN_815;
  assign _GEN_880 = 6'he == _T_218 ? _GEN_13 : _GEN_816;
  assign _GEN_881 = 6'hf == _T_218 ? _GEN_13 : _GEN_817;
  assign _GEN_882 = 6'h10 == _T_218 ? _GEN_13 : _GEN_818;
  assign _GEN_883 = 6'h11 == _T_218 ? _GEN_13 : _GEN_819;
  assign _GEN_884 = 6'h12 == _T_218 ? _GEN_13 : _GEN_820;
  assign _GEN_885 = 6'h13 == _T_218 ? _GEN_13 : _GEN_821;
  assign _GEN_886 = 6'h14 == _T_218 ? _GEN_13 : _GEN_822;
  assign _GEN_887 = 6'h15 == _T_218 ? _GEN_13 : _GEN_823;
  assign _GEN_888 = 6'h16 == _T_218 ? _GEN_13 : _GEN_824;
  assign _GEN_889 = 6'h17 == _T_218 ? _GEN_13 : _GEN_825;
  assign _GEN_890 = 6'h18 == _T_218 ? _GEN_13 : _GEN_826;
  assign _GEN_891 = 6'h19 == _T_218 ? _GEN_13 : _GEN_827;
  assign _GEN_892 = 6'h1a == _T_218 ? _GEN_13 : _GEN_828;
  assign _GEN_893 = 6'h1b == _T_218 ? _GEN_13 : _GEN_829;
  assign _GEN_894 = 6'h1c == _T_218 ? _GEN_13 : _GEN_830;
  assign _GEN_895 = 6'h1d == _T_218 ? _GEN_13 : _GEN_831;
  assign _GEN_896 = 6'h1e == _T_218 ? _GEN_13 : _GEN_832;
  assign _GEN_897 = 6'h1f == _T_218 ? _GEN_13 : _GEN_833;
  assign _GEN_898 = 6'h20 == _T_218 ? _GEN_13 : _GEN_834;
  assign _GEN_899 = 6'h21 == _T_218 ? _GEN_13 : _GEN_835;
  assign _GEN_900 = 6'h22 == _T_218 ? _GEN_13 : _GEN_836;
  assign _GEN_901 = 6'h23 == _T_218 ? _GEN_13 : _GEN_837;
  assign _GEN_902 = 6'h24 == _T_218 ? _GEN_13 : _GEN_838;
  assign _GEN_903 = 6'h25 == _T_218 ? _GEN_13 : _GEN_839;
  assign _GEN_904 = 6'h26 == _T_218 ? _GEN_13 : _GEN_840;
  assign _GEN_905 = 6'h27 == _T_218 ? _GEN_13 : _GEN_841;
  assign _GEN_906 = 6'h28 == _T_218 ? _GEN_13 : _GEN_842;
  assign _GEN_907 = 6'h29 == _T_218 ? _GEN_13 : _GEN_843;
  assign _GEN_908 = 6'h2a == _T_218 ? _GEN_13 : _GEN_844;
  assign _GEN_909 = 6'h2b == _T_218 ? _GEN_13 : _GEN_845;
  assign _GEN_910 = 6'h2c == _T_218 ? _GEN_13 : _GEN_846;
  assign _GEN_911 = 6'h2d == _T_218 ? _GEN_13 : _GEN_847;
  assign _GEN_912 = 6'h2e == _T_218 ? _GEN_13 : _GEN_848;
  assign _GEN_913 = 6'h2f == _T_218 ? _GEN_13 : _GEN_849;
  assign _GEN_914 = 6'h30 == _T_218 ? _GEN_13 : _GEN_850;
  assign _GEN_915 = 6'h31 == _T_218 ? _GEN_13 : _GEN_851;
  assign _GEN_916 = 6'h32 == _T_218 ? _GEN_13 : _GEN_852;
  assign _GEN_917 = 6'h33 == _T_218 ? _GEN_13 : _GEN_853;
  assign _GEN_918 = 6'h34 == _T_218 ? _GEN_13 : _GEN_854;
  assign _GEN_919 = 6'h35 == _T_218 ? _GEN_13 : _GEN_855;
  assign _GEN_920 = 6'h36 == _T_218 ? _GEN_13 : _GEN_856;
  assign _GEN_921 = 6'h37 == _T_218 ? _GEN_13 : _GEN_857;
  assign _GEN_922 = 6'h38 == _T_218 ? _GEN_13 : _GEN_858;
  assign _GEN_923 = 6'h39 == _T_218 ? _GEN_13 : _GEN_859;
  assign _GEN_924 = 6'h3a == _T_218 ? _GEN_13 : _GEN_860;
  assign _GEN_925 = 6'h3b == _T_218 ? _GEN_13 : _GEN_861;
  assign _GEN_926 = 6'h3c == _T_218 ? _GEN_13 : _GEN_862;
  assign _GEN_927 = 6'h3d == _T_218 ? _GEN_13 : _GEN_863;
  assign _GEN_928 = 6'h3e == _T_218 ? _GEN_13 : _GEN_864;
  assign _GEN_929 = 6'h3f == _T_218 ? _GEN_13 : _GEN_865;
  assign _T_222 = wPos + 6'he;
  assign _T_223 = _T_222[5:0];
  assign _T_225 = io_fastin[71:68];
  assign _GEN_14 = _T_225;
  assign _GEN_930 = 6'h0 == _T_223 ? _GEN_14 : _GEN_866;
  assign _GEN_931 = 6'h1 == _T_223 ? _GEN_14 : _GEN_867;
  assign _GEN_932 = 6'h2 == _T_223 ? _GEN_14 : _GEN_868;
  assign _GEN_933 = 6'h3 == _T_223 ? _GEN_14 : _GEN_869;
  assign _GEN_934 = 6'h4 == _T_223 ? _GEN_14 : _GEN_870;
  assign _GEN_935 = 6'h5 == _T_223 ? _GEN_14 : _GEN_871;
  assign _GEN_936 = 6'h6 == _T_223 ? _GEN_14 : _GEN_872;
  assign _GEN_937 = 6'h7 == _T_223 ? _GEN_14 : _GEN_873;
  assign _GEN_938 = 6'h8 == _T_223 ? _GEN_14 : _GEN_874;
  assign _GEN_939 = 6'h9 == _T_223 ? _GEN_14 : _GEN_875;
  assign _GEN_940 = 6'ha == _T_223 ? _GEN_14 : _GEN_876;
  assign _GEN_941 = 6'hb == _T_223 ? _GEN_14 : _GEN_877;
  assign _GEN_942 = 6'hc == _T_223 ? _GEN_14 : _GEN_878;
  assign _GEN_943 = 6'hd == _T_223 ? _GEN_14 : _GEN_879;
  assign _GEN_944 = 6'he == _T_223 ? _GEN_14 : _GEN_880;
  assign _GEN_945 = 6'hf == _T_223 ? _GEN_14 : _GEN_881;
  assign _GEN_946 = 6'h10 == _T_223 ? _GEN_14 : _GEN_882;
  assign _GEN_947 = 6'h11 == _T_223 ? _GEN_14 : _GEN_883;
  assign _GEN_948 = 6'h12 == _T_223 ? _GEN_14 : _GEN_884;
  assign _GEN_949 = 6'h13 == _T_223 ? _GEN_14 : _GEN_885;
  assign _GEN_950 = 6'h14 == _T_223 ? _GEN_14 : _GEN_886;
  assign _GEN_951 = 6'h15 == _T_223 ? _GEN_14 : _GEN_887;
  assign _GEN_952 = 6'h16 == _T_223 ? _GEN_14 : _GEN_888;
  assign _GEN_953 = 6'h17 == _T_223 ? _GEN_14 : _GEN_889;
  assign _GEN_954 = 6'h18 == _T_223 ? _GEN_14 : _GEN_890;
  assign _GEN_955 = 6'h19 == _T_223 ? _GEN_14 : _GEN_891;
  assign _GEN_956 = 6'h1a == _T_223 ? _GEN_14 : _GEN_892;
  assign _GEN_957 = 6'h1b == _T_223 ? _GEN_14 : _GEN_893;
  assign _GEN_958 = 6'h1c == _T_223 ? _GEN_14 : _GEN_894;
  assign _GEN_959 = 6'h1d == _T_223 ? _GEN_14 : _GEN_895;
  assign _GEN_960 = 6'h1e == _T_223 ? _GEN_14 : _GEN_896;
  assign _GEN_961 = 6'h1f == _T_223 ? _GEN_14 : _GEN_897;
  assign _GEN_962 = 6'h20 == _T_223 ? _GEN_14 : _GEN_898;
  assign _GEN_963 = 6'h21 == _T_223 ? _GEN_14 : _GEN_899;
  assign _GEN_964 = 6'h22 == _T_223 ? _GEN_14 : _GEN_900;
  assign _GEN_965 = 6'h23 == _T_223 ? _GEN_14 : _GEN_901;
  assign _GEN_966 = 6'h24 == _T_223 ? _GEN_14 : _GEN_902;
  assign _GEN_967 = 6'h25 == _T_223 ? _GEN_14 : _GEN_903;
  assign _GEN_968 = 6'h26 == _T_223 ? _GEN_14 : _GEN_904;
  assign _GEN_969 = 6'h27 == _T_223 ? _GEN_14 : _GEN_905;
  assign _GEN_970 = 6'h28 == _T_223 ? _GEN_14 : _GEN_906;
  assign _GEN_971 = 6'h29 == _T_223 ? _GEN_14 : _GEN_907;
  assign _GEN_972 = 6'h2a == _T_223 ? _GEN_14 : _GEN_908;
  assign _GEN_973 = 6'h2b == _T_223 ? _GEN_14 : _GEN_909;
  assign _GEN_974 = 6'h2c == _T_223 ? _GEN_14 : _GEN_910;
  assign _GEN_975 = 6'h2d == _T_223 ? _GEN_14 : _GEN_911;
  assign _GEN_976 = 6'h2e == _T_223 ? _GEN_14 : _GEN_912;
  assign _GEN_977 = 6'h2f == _T_223 ? _GEN_14 : _GEN_913;
  assign _GEN_978 = 6'h30 == _T_223 ? _GEN_14 : _GEN_914;
  assign _GEN_979 = 6'h31 == _T_223 ? _GEN_14 : _GEN_915;
  assign _GEN_980 = 6'h32 == _T_223 ? _GEN_14 : _GEN_916;
  assign _GEN_981 = 6'h33 == _T_223 ? _GEN_14 : _GEN_917;
  assign _GEN_982 = 6'h34 == _T_223 ? _GEN_14 : _GEN_918;
  assign _GEN_983 = 6'h35 == _T_223 ? _GEN_14 : _GEN_919;
  assign _GEN_984 = 6'h36 == _T_223 ? _GEN_14 : _GEN_920;
  assign _GEN_985 = 6'h37 == _T_223 ? _GEN_14 : _GEN_921;
  assign _GEN_986 = 6'h38 == _T_223 ? _GEN_14 : _GEN_922;
  assign _GEN_987 = 6'h39 == _T_223 ? _GEN_14 : _GEN_923;
  assign _GEN_988 = 6'h3a == _T_223 ? _GEN_14 : _GEN_924;
  assign _GEN_989 = 6'h3b == _T_223 ? _GEN_14 : _GEN_925;
  assign _GEN_990 = 6'h3c == _T_223 ? _GEN_14 : _GEN_926;
  assign _GEN_991 = 6'h3d == _T_223 ? _GEN_14 : _GEN_927;
  assign _GEN_992 = 6'h3e == _T_223 ? _GEN_14 : _GEN_928;
  assign _GEN_993 = 6'h3f == _T_223 ? _GEN_14 : _GEN_929;
  assign _T_227 = wPos + 6'hf;
  assign _T_228 = _T_227[5:0];
  assign _T_230 = io_fastin[67:64];
  assign _GEN_15 = _T_230;
  assign _GEN_994 = 6'h0 == _T_228 ? _GEN_15 : _GEN_930;
  assign _GEN_995 = 6'h1 == _T_228 ? _GEN_15 : _GEN_931;
  assign _GEN_996 = 6'h2 == _T_228 ? _GEN_15 : _GEN_932;
  assign _GEN_997 = 6'h3 == _T_228 ? _GEN_15 : _GEN_933;
  assign _GEN_998 = 6'h4 == _T_228 ? _GEN_15 : _GEN_934;
  assign _GEN_999 = 6'h5 == _T_228 ? _GEN_15 : _GEN_935;
  assign _GEN_1000 = 6'h6 == _T_228 ? _GEN_15 : _GEN_936;
  assign _GEN_1001 = 6'h7 == _T_228 ? _GEN_15 : _GEN_937;
  assign _GEN_1002 = 6'h8 == _T_228 ? _GEN_15 : _GEN_938;
  assign _GEN_1003 = 6'h9 == _T_228 ? _GEN_15 : _GEN_939;
  assign _GEN_1004 = 6'ha == _T_228 ? _GEN_15 : _GEN_940;
  assign _GEN_1005 = 6'hb == _T_228 ? _GEN_15 : _GEN_941;
  assign _GEN_1006 = 6'hc == _T_228 ? _GEN_15 : _GEN_942;
  assign _GEN_1007 = 6'hd == _T_228 ? _GEN_15 : _GEN_943;
  assign _GEN_1008 = 6'he == _T_228 ? _GEN_15 : _GEN_944;
  assign _GEN_1009 = 6'hf == _T_228 ? _GEN_15 : _GEN_945;
  assign _GEN_1010 = 6'h10 == _T_228 ? _GEN_15 : _GEN_946;
  assign _GEN_1011 = 6'h11 == _T_228 ? _GEN_15 : _GEN_947;
  assign _GEN_1012 = 6'h12 == _T_228 ? _GEN_15 : _GEN_948;
  assign _GEN_1013 = 6'h13 == _T_228 ? _GEN_15 : _GEN_949;
  assign _GEN_1014 = 6'h14 == _T_228 ? _GEN_15 : _GEN_950;
  assign _GEN_1015 = 6'h15 == _T_228 ? _GEN_15 : _GEN_951;
  assign _GEN_1016 = 6'h16 == _T_228 ? _GEN_15 : _GEN_952;
  assign _GEN_1017 = 6'h17 == _T_228 ? _GEN_15 : _GEN_953;
  assign _GEN_1018 = 6'h18 == _T_228 ? _GEN_15 : _GEN_954;
  assign _GEN_1019 = 6'h19 == _T_228 ? _GEN_15 : _GEN_955;
  assign _GEN_1020 = 6'h1a == _T_228 ? _GEN_15 : _GEN_956;
  assign _GEN_1021 = 6'h1b == _T_228 ? _GEN_15 : _GEN_957;
  assign _GEN_1022 = 6'h1c == _T_228 ? _GEN_15 : _GEN_958;
  assign _GEN_1023 = 6'h1d == _T_228 ? _GEN_15 : _GEN_959;
  assign _GEN_1024 = 6'h1e == _T_228 ? _GEN_15 : _GEN_960;
  assign _GEN_1025 = 6'h1f == _T_228 ? _GEN_15 : _GEN_961;
  assign _GEN_1026 = 6'h20 == _T_228 ? _GEN_15 : _GEN_962;
  assign _GEN_1027 = 6'h21 == _T_228 ? _GEN_15 : _GEN_963;
  assign _GEN_1028 = 6'h22 == _T_228 ? _GEN_15 : _GEN_964;
  assign _GEN_1029 = 6'h23 == _T_228 ? _GEN_15 : _GEN_965;
  assign _GEN_1030 = 6'h24 == _T_228 ? _GEN_15 : _GEN_966;
  assign _GEN_1031 = 6'h25 == _T_228 ? _GEN_15 : _GEN_967;
  assign _GEN_1032 = 6'h26 == _T_228 ? _GEN_15 : _GEN_968;
  assign _GEN_1033 = 6'h27 == _T_228 ? _GEN_15 : _GEN_969;
  assign _GEN_1034 = 6'h28 == _T_228 ? _GEN_15 : _GEN_970;
  assign _GEN_1035 = 6'h29 == _T_228 ? _GEN_15 : _GEN_971;
  assign _GEN_1036 = 6'h2a == _T_228 ? _GEN_15 : _GEN_972;
  assign _GEN_1037 = 6'h2b == _T_228 ? _GEN_15 : _GEN_973;
  assign _GEN_1038 = 6'h2c == _T_228 ? _GEN_15 : _GEN_974;
  assign _GEN_1039 = 6'h2d == _T_228 ? _GEN_15 : _GEN_975;
  assign _GEN_1040 = 6'h2e == _T_228 ? _GEN_15 : _GEN_976;
  assign _GEN_1041 = 6'h2f == _T_228 ? _GEN_15 : _GEN_977;
  assign _GEN_1042 = 6'h30 == _T_228 ? _GEN_15 : _GEN_978;
  assign _GEN_1043 = 6'h31 == _T_228 ? _GEN_15 : _GEN_979;
  assign _GEN_1044 = 6'h32 == _T_228 ? _GEN_15 : _GEN_980;
  assign _GEN_1045 = 6'h33 == _T_228 ? _GEN_15 : _GEN_981;
  assign _GEN_1046 = 6'h34 == _T_228 ? _GEN_15 : _GEN_982;
  assign _GEN_1047 = 6'h35 == _T_228 ? _GEN_15 : _GEN_983;
  assign _GEN_1048 = 6'h36 == _T_228 ? _GEN_15 : _GEN_984;
  assign _GEN_1049 = 6'h37 == _T_228 ? _GEN_15 : _GEN_985;
  assign _GEN_1050 = 6'h38 == _T_228 ? _GEN_15 : _GEN_986;
  assign _GEN_1051 = 6'h39 == _T_228 ? _GEN_15 : _GEN_987;
  assign _GEN_1052 = 6'h3a == _T_228 ? _GEN_15 : _GEN_988;
  assign _GEN_1053 = 6'h3b == _T_228 ? _GEN_15 : _GEN_989;
  assign _GEN_1054 = 6'h3c == _T_228 ? _GEN_15 : _GEN_990;
  assign _GEN_1055 = 6'h3d == _T_228 ? _GEN_15 : _GEN_991;
  assign _GEN_1056 = 6'h3e == _T_228 ? _GEN_15 : _GEN_992;
  assign _GEN_1057 = 6'h3f == _T_228 ? _GEN_15 : _GEN_993;
  assign _T_232 = wPos + 6'h10;
  assign _T_233 = _T_232[5:0];
  assign _T_235 = io_fastin[63:60];
  assign _GEN_16 = _T_235;
  assign _GEN_1058 = 6'h0 == _T_233 ? _GEN_16 : _GEN_994;
  assign _GEN_1059 = 6'h1 == _T_233 ? _GEN_16 : _GEN_995;
  assign _GEN_1060 = 6'h2 == _T_233 ? _GEN_16 : _GEN_996;
  assign _GEN_1061 = 6'h3 == _T_233 ? _GEN_16 : _GEN_997;
  assign _GEN_1062 = 6'h4 == _T_233 ? _GEN_16 : _GEN_998;
  assign _GEN_1063 = 6'h5 == _T_233 ? _GEN_16 : _GEN_999;
  assign _GEN_1064 = 6'h6 == _T_233 ? _GEN_16 : _GEN_1000;
  assign _GEN_1065 = 6'h7 == _T_233 ? _GEN_16 : _GEN_1001;
  assign _GEN_1066 = 6'h8 == _T_233 ? _GEN_16 : _GEN_1002;
  assign _GEN_1067 = 6'h9 == _T_233 ? _GEN_16 : _GEN_1003;
  assign _GEN_1068 = 6'ha == _T_233 ? _GEN_16 : _GEN_1004;
  assign _GEN_1069 = 6'hb == _T_233 ? _GEN_16 : _GEN_1005;
  assign _GEN_1070 = 6'hc == _T_233 ? _GEN_16 : _GEN_1006;
  assign _GEN_1071 = 6'hd == _T_233 ? _GEN_16 : _GEN_1007;
  assign _GEN_1072 = 6'he == _T_233 ? _GEN_16 : _GEN_1008;
  assign _GEN_1073 = 6'hf == _T_233 ? _GEN_16 : _GEN_1009;
  assign _GEN_1074 = 6'h10 == _T_233 ? _GEN_16 : _GEN_1010;
  assign _GEN_1075 = 6'h11 == _T_233 ? _GEN_16 : _GEN_1011;
  assign _GEN_1076 = 6'h12 == _T_233 ? _GEN_16 : _GEN_1012;
  assign _GEN_1077 = 6'h13 == _T_233 ? _GEN_16 : _GEN_1013;
  assign _GEN_1078 = 6'h14 == _T_233 ? _GEN_16 : _GEN_1014;
  assign _GEN_1079 = 6'h15 == _T_233 ? _GEN_16 : _GEN_1015;
  assign _GEN_1080 = 6'h16 == _T_233 ? _GEN_16 : _GEN_1016;
  assign _GEN_1081 = 6'h17 == _T_233 ? _GEN_16 : _GEN_1017;
  assign _GEN_1082 = 6'h18 == _T_233 ? _GEN_16 : _GEN_1018;
  assign _GEN_1083 = 6'h19 == _T_233 ? _GEN_16 : _GEN_1019;
  assign _GEN_1084 = 6'h1a == _T_233 ? _GEN_16 : _GEN_1020;
  assign _GEN_1085 = 6'h1b == _T_233 ? _GEN_16 : _GEN_1021;
  assign _GEN_1086 = 6'h1c == _T_233 ? _GEN_16 : _GEN_1022;
  assign _GEN_1087 = 6'h1d == _T_233 ? _GEN_16 : _GEN_1023;
  assign _GEN_1088 = 6'h1e == _T_233 ? _GEN_16 : _GEN_1024;
  assign _GEN_1089 = 6'h1f == _T_233 ? _GEN_16 : _GEN_1025;
  assign _GEN_1090 = 6'h20 == _T_233 ? _GEN_16 : _GEN_1026;
  assign _GEN_1091 = 6'h21 == _T_233 ? _GEN_16 : _GEN_1027;
  assign _GEN_1092 = 6'h22 == _T_233 ? _GEN_16 : _GEN_1028;
  assign _GEN_1093 = 6'h23 == _T_233 ? _GEN_16 : _GEN_1029;
  assign _GEN_1094 = 6'h24 == _T_233 ? _GEN_16 : _GEN_1030;
  assign _GEN_1095 = 6'h25 == _T_233 ? _GEN_16 : _GEN_1031;
  assign _GEN_1096 = 6'h26 == _T_233 ? _GEN_16 : _GEN_1032;
  assign _GEN_1097 = 6'h27 == _T_233 ? _GEN_16 : _GEN_1033;
  assign _GEN_1098 = 6'h28 == _T_233 ? _GEN_16 : _GEN_1034;
  assign _GEN_1099 = 6'h29 == _T_233 ? _GEN_16 : _GEN_1035;
  assign _GEN_1100 = 6'h2a == _T_233 ? _GEN_16 : _GEN_1036;
  assign _GEN_1101 = 6'h2b == _T_233 ? _GEN_16 : _GEN_1037;
  assign _GEN_1102 = 6'h2c == _T_233 ? _GEN_16 : _GEN_1038;
  assign _GEN_1103 = 6'h2d == _T_233 ? _GEN_16 : _GEN_1039;
  assign _GEN_1104 = 6'h2e == _T_233 ? _GEN_16 : _GEN_1040;
  assign _GEN_1105 = 6'h2f == _T_233 ? _GEN_16 : _GEN_1041;
  assign _GEN_1106 = 6'h30 == _T_233 ? _GEN_16 : _GEN_1042;
  assign _GEN_1107 = 6'h31 == _T_233 ? _GEN_16 : _GEN_1043;
  assign _GEN_1108 = 6'h32 == _T_233 ? _GEN_16 : _GEN_1044;
  assign _GEN_1109 = 6'h33 == _T_233 ? _GEN_16 : _GEN_1045;
  assign _GEN_1110 = 6'h34 == _T_233 ? _GEN_16 : _GEN_1046;
  assign _GEN_1111 = 6'h35 == _T_233 ? _GEN_16 : _GEN_1047;
  assign _GEN_1112 = 6'h36 == _T_233 ? _GEN_16 : _GEN_1048;
  assign _GEN_1113 = 6'h37 == _T_233 ? _GEN_16 : _GEN_1049;
  assign _GEN_1114 = 6'h38 == _T_233 ? _GEN_16 : _GEN_1050;
  assign _GEN_1115 = 6'h39 == _T_233 ? _GEN_16 : _GEN_1051;
  assign _GEN_1116 = 6'h3a == _T_233 ? _GEN_16 : _GEN_1052;
  assign _GEN_1117 = 6'h3b == _T_233 ? _GEN_16 : _GEN_1053;
  assign _GEN_1118 = 6'h3c == _T_233 ? _GEN_16 : _GEN_1054;
  assign _GEN_1119 = 6'h3d == _T_233 ? _GEN_16 : _GEN_1055;
  assign _GEN_1120 = 6'h3e == _T_233 ? _GEN_16 : _GEN_1056;
  assign _GEN_1121 = 6'h3f == _T_233 ? _GEN_16 : _GEN_1057;
  assign _T_237 = wPos + 6'h11;
  assign _T_238 = _T_237[5:0];
  assign _T_240 = io_fastin[59:56];
  assign _GEN_17 = _T_240;
  assign _GEN_1122 = 6'h0 == _T_238 ? _GEN_17 : _GEN_1058;
  assign _GEN_1123 = 6'h1 == _T_238 ? _GEN_17 : _GEN_1059;
  assign _GEN_1124 = 6'h2 == _T_238 ? _GEN_17 : _GEN_1060;
  assign _GEN_1125 = 6'h3 == _T_238 ? _GEN_17 : _GEN_1061;
  assign _GEN_1126 = 6'h4 == _T_238 ? _GEN_17 : _GEN_1062;
  assign _GEN_1127 = 6'h5 == _T_238 ? _GEN_17 : _GEN_1063;
  assign _GEN_1128 = 6'h6 == _T_238 ? _GEN_17 : _GEN_1064;
  assign _GEN_1129 = 6'h7 == _T_238 ? _GEN_17 : _GEN_1065;
  assign _GEN_1130 = 6'h8 == _T_238 ? _GEN_17 : _GEN_1066;
  assign _GEN_1131 = 6'h9 == _T_238 ? _GEN_17 : _GEN_1067;
  assign _GEN_1132 = 6'ha == _T_238 ? _GEN_17 : _GEN_1068;
  assign _GEN_1133 = 6'hb == _T_238 ? _GEN_17 : _GEN_1069;
  assign _GEN_1134 = 6'hc == _T_238 ? _GEN_17 : _GEN_1070;
  assign _GEN_1135 = 6'hd == _T_238 ? _GEN_17 : _GEN_1071;
  assign _GEN_1136 = 6'he == _T_238 ? _GEN_17 : _GEN_1072;
  assign _GEN_1137 = 6'hf == _T_238 ? _GEN_17 : _GEN_1073;
  assign _GEN_1138 = 6'h10 == _T_238 ? _GEN_17 : _GEN_1074;
  assign _GEN_1139 = 6'h11 == _T_238 ? _GEN_17 : _GEN_1075;
  assign _GEN_1140 = 6'h12 == _T_238 ? _GEN_17 : _GEN_1076;
  assign _GEN_1141 = 6'h13 == _T_238 ? _GEN_17 : _GEN_1077;
  assign _GEN_1142 = 6'h14 == _T_238 ? _GEN_17 : _GEN_1078;
  assign _GEN_1143 = 6'h15 == _T_238 ? _GEN_17 : _GEN_1079;
  assign _GEN_1144 = 6'h16 == _T_238 ? _GEN_17 : _GEN_1080;
  assign _GEN_1145 = 6'h17 == _T_238 ? _GEN_17 : _GEN_1081;
  assign _GEN_1146 = 6'h18 == _T_238 ? _GEN_17 : _GEN_1082;
  assign _GEN_1147 = 6'h19 == _T_238 ? _GEN_17 : _GEN_1083;
  assign _GEN_1148 = 6'h1a == _T_238 ? _GEN_17 : _GEN_1084;
  assign _GEN_1149 = 6'h1b == _T_238 ? _GEN_17 : _GEN_1085;
  assign _GEN_1150 = 6'h1c == _T_238 ? _GEN_17 : _GEN_1086;
  assign _GEN_1151 = 6'h1d == _T_238 ? _GEN_17 : _GEN_1087;
  assign _GEN_1152 = 6'h1e == _T_238 ? _GEN_17 : _GEN_1088;
  assign _GEN_1153 = 6'h1f == _T_238 ? _GEN_17 : _GEN_1089;
  assign _GEN_1154 = 6'h20 == _T_238 ? _GEN_17 : _GEN_1090;
  assign _GEN_1155 = 6'h21 == _T_238 ? _GEN_17 : _GEN_1091;
  assign _GEN_1156 = 6'h22 == _T_238 ? _GEN_17 : _GEN_1092;
  assign _GEN_1157 = 6'h23 == _T_238 ? _GEN_17 : _GEN_1093;
  assign _GEN_1158 = 6'h24 == _T_238 ? _GEN_17 : _GEN_1094;
  assign _GEN_1159 = 6'h25 == _T_238 ? _GEN_17 : _GEN_1095;
  assign _GEN_1160 = 6'h26 == _T_238 ? _GEN_17 : _GEN_1096;
  assign _GEN_1161 = 6'h27 == _T_238 ? _GEN_17 : _GEN_1097;
  assign _GEN_1162 = 6'h28 == _T_238 ? _GEN_17 : _GEN_1098;
  assign _GEN_1163 = 6'h29 == _T_238 ? _GEN_17 : _GEN_1099;
  assign _GEN_1164 = 6'h2a == _T_238 ? _GEN_17 : _GEN_1100;
  assign _GEN_1165 = 6'h2b == _T_238 ? _GEN_17 : _GEN_1101;
  assign _GEN_1166 = 6'h2c == _T_238 ? _GEN_17 : _GEN_1102;
  assign _GEN_1167 = 6'h2d == _T_238 ? _GEN_17 : _GEN_1103;
  assign _GEN_1168 = 6'h2e == _T_238 ? _GEN_17 : _GEN_1104;
  assign _GEN_1169 = 6'h2f == _T_238 ? _GEN_17 : _GEN_1105;
  assign _GEN_1170 = 6'h30 == _T_238 ? _GEN_17 : _GEN_1106;
  assign _GEN_1171 = 6'h31 == _T_238 ? _GEN_17 : _GEN_1107;
  assign _GEN_1172 = 6'h32 == _T_238 ? _GEN_17 : _GEN_1108;
  assign _GEN_1173 = 6'h33 == _T_238 ? _GEN_17 : _GEN_1109;
  assign _GEN_1174 = 6'h34 == _T_238 ? _GEN_17 : _GEN_1110;
  assign _GEN_1175 = 6'h35 == _T_238 ? _GEN_17 : _GEN_1111;
  assign _GEN_1176 = 6'h36 == _T_238 ? _GEN_17 : _GEN_1112;
  assign _GEN_1177 = 6'h37 == _T_238 ? _GEN_17 : _GEN_1113;
  assign _GEN_1178 = 6'h38 == _T_238 ? _GEN_17 : _GEN_1114;
  assign _GEN_1179 = 6'h39 == _T_238 ? _GEN_17 : _GEN_1115;
  assign _GEN_1180 = 6'h3a == _T_238 ? _GEN_17 : _GEN_1116;
  assign _GEN_1181 = 6'h3b == _T_238 ? _GEN_17 : _GEN_1117;
  assign _GEN_1182 = 6'h3c == _T_238 ? _GEN_17 : _GEN_1118;
  assign _GEN_1183 = 6'h3d == _T_238 ? _GEN_17 : _GEN_1119;
  assign _GEN_1184 = 6'h3e == _T_238 ? _GEN_17 : _GEN_1120;
  assign _GEN_1185 = 6'h3f == _T_238 ? _GEN_17 : _GEN_1121;
  assign _T_242 = wPos + 6'h12;
  assign _T_243 = _T_242[5:0];
  assign _T_245 = io_fastin[55:52];
  assign _GEN_18 = _T_245;
  assign _GEN_1186 = 6'h0 == _T_243 ? _GEN_18 : _GEN_1122;
  assign _GEN_1187 = 6'h1 == _T_243 ? _GEN_18 : _GEN_1123;
  assign _GEN_1188 = 6'h2 == _T_243 ? _GEN_18 : _GEN_1124;
  assign _GEN_1189 = 6'h3 == _T_243 ? _GEN_18 : _GEN_1125;
  assign _GEN_1190 = 6'h4 == _T_243 ? _GEN_18 : _GEN_1126;
  assign _GEN_1191 = 6'h5 == _T_243 ? _GEN_18 : _GEN_1127;
  assign _GEN_1192 = 6'h6 == _T_243 ? _GEN_18 : _GEN_1128;
  assign _GEN_1193 = 6'h7 == _T_243 ? _GEN_18 : _GEN_1129;
  assign _GEN_1194 = 6'h8 == _T_243 ? _GEN_18 : _GEN_1130;
  assign _GEN_1195 = 6'h9 == _T_243 ? _GEN_18 : _GEN_1131;
  assign _GEN_1196 = 6'ha == _T_243 ? _GEN_18 : _GEN_1132;
  assign _GEN_1197 = 6'hb == _T_243 ? _GEN_18 : _GEN_1133;
  assign _GEN_1198 = 6'hc == _T_243 ? _GEN_18 : _GEN_1134;
  assign _GEN_1199 = 6'hd == _T_243 ? _GEN_18 : _GEN_1135;
  assign _GEN_1200 = 6'he == _T_243 ? _GEN_18 : _GEN_1136;
  assign _GEN_1201 = 6'hf == _T_243 ? _GEN_18 : _GEN_1137;
  assign _GEN_1202 = 6'h10 == _T_243 ? _GEN_18 : _GEN_1138;
  assign _GEN_1203 = 6'h11 == _T_243 ? _GEN_18 : _GEN_1139;
  assign _GEN_1204 = 6'h12 == _T_243 ? _GEN_18 : _GEN_1140;
  assign _GEN_1205 = 6'h13 == _T_243 ? _GEN_18 : _GEN_1141;
  assign _GEN_1206 = 6'h14 == _T_243 ? _GEN_18 : _GEN_1142;
  assign _GEN_1207 = 6'h15 == _T_243 ? _GEN_18 : _GEN_1143;
  assign _GEN_1208 = 6'h16 == _T_243 ? _GEN_18 : _GEN_1144;
  assign _GEN_1209 = 6'h17 == _T_243 ? _GEN_18 : _GEN_1145;
  assign _GEN_1210 = 6'h18 == _T_243 ? _GEN_18 : _GEN_1146;
  assign _GEN_1211 = 6'h19 == _T_243 ? _GEN_18 : _GEN_1147;
  assign _GEN_1212 = 6'h1a == _T_243 ? _GEN_18 : _GEN_1148;
  assign _GEN_1213 = 6'h1b == _T_243 ? _GEN_18 : _GEN_1149;
  assign _GEN_1214 = 6'h1c == _T_243 ? _GEN_18 : _GEN_1150;
  assign _GEN_1215 = 6'h1d == _T_243 ? _GEN_18 : _GEN_1151;
  assign _GEN_1216 = 6'h1e == _T_243 ? _GEN_18 : _GEN_1152;
  assign _GEN_1217 = 6'h1f == _T_243 ? _GEN_18 : _GEN_1153;
  assign _GEN_1218 = 6'h20 == _T_243 ? _GEN_18 : _GEN_1154;
  assign _GEN_1219 = 6'h21 == _T_243 ? _GEN_18 : _GEN_1155;
  assign _GEN_1220 = 6'h22 == _T_243 ? _GEN_18 : _GEN_1156;
  assign _GEN_1221 = 6'h23 == _T_243 ? _GEN_18 : _GEN_1157;
  assign _GEN_1222 = 6'h24 == _T_243 ? _GEN_18 : _GEN_1158;
  assign _GEN_1223 = 6'h25 == _T_243 ? _GEN_18 : _GEN_1159;
  assign _GEN_1224 = 6'h26 == _T_243 ? _GEN_18 : _GEN_1160;
  assign _GEN_1225 = 6'h27 == _T_243 ? _GEN_18 : _GEN_1161;
  assign _GEN_1226 = 6'h28 == _T_243 ? _GEN_18 : _GEN_1162;
  assign _GEN_1227 = 6'h29 == _T_243 ? _GEN_18 : _GEN_1163;
  assign _GEN_1228 = 6'h2a == _T_243 ? _GEN_18 : _GEN_1164;
  assign _GEN_1229 = 6'h2b == _T_243 ? _GEN_18 : _GEN_1165;
  assign _GEN_1230 = 6'h2c == _T_243 ? _GEN_18 : _GEN_1166;
  assign _GEN_1231 = 6'h2d == _T_243 ? _GEN_18 : _GEN_1167;
  assign _GEN_1232 = 6'h2e == _T_243 ? _GEN_18 : _GEN_1168;
  assign _GEN_1233 = 6'h2f == _T_243 ? _GEN_18 : _GEN_1169;
  assign _GEN_1234 = 6'h30 == _T_243 ? _GEN_18 : _GEN_1170;
  assign _GEN_1235 = 6'h31 == _T_243 ? _GEN_18 : _GEN_1171;
  assign _GEN_1236 = 6'h32 == _T_243 ? _GEN_18 : _GEN_1172;
  assign _GEN_1237 = 6'h33 == _T_243 ? _GEN_18 : _GEN_1173;
  assign _GEN_1238 = 6'h34 == _T_243 ? _GEN_18 : _GEN_1174;
  assign _GEN_1239 = 6'h35 == _T_243 ? _GEN_18 : _GEN_1175;
  assign _GEN_1240 = 6'h36 == _T_243 ? _GEN_18 : _GEN_1176;
  assign _GEN_1241 = 6'h37 == _T_243 ? _GEN_18 : _GEN_1177;
  assign _GEN_1242 = 6'h38 == _T_243 ? _GEN_18 : _GEN_1178;
  assign _GEN_1243 = 6'h39 == _T_243 ? _GEN_18 : _GEN_1179;
  assign _GEN_1244 = 6'h3a == _T_243 ? _GEN_18 : _GEN_1180;
  assign _GEN_1245 = 6'h3b == _T_243 ? _GEN_18 : _GEN_1181;
  assign _GEN_1246 = 6'h3c == _T_243 ? _GEN_18 : _GEN_1182;
  assign _GEN_1247 = 6'h3d == _T_243 ? _GEN_18 : _GEN_1183;
  assign _GEN_1248 = 6'h3e == _T_243 ? _GEN_18 : _GEN_1184;
  assign _GEN_1249 = 6'h3f == _T_243 ? _GEN_18 : _GEN_1185;
  assign _T_247 = wPos + 6'h13;
  assign _T_248 = _T_247[5:0];
  assign _T_250 = io_fastin[51:48];
  assign _GEN_19 = _T_250;
  assign _GEN_1250 = 6'h0 == _T_248 ? _GEN_19 : _GEN_1186;
  assign _GEN_1251 = 6'h1 == _T_248 ? _GEN_19 : _GEN_1187;
  assign _GEN_1252 = 6'h2 == _T_248 ? _GEN_19 : _GEN_1188;
  assign _GEN_1253 = 6'h3 == _T_248 ? _GEN_19 : _GEN_1189;
  assign _GEN_1254 = 6'h4 == _T_248 ? _GEN_19 : _GEN_1190;
  assign _GEN_1255 = 6'h5 == _T_248 ? _GEN_19 : _GEN_1191;
  assign _GEN_1256 = 6'h6 == _T_248 ? _GEN_19 : _GEN_1192;
  assign _GEN_1257 = 6'h7 == _T_248 ? _GEN_19 : _GEN_1193;
  assign _GEN_1258 = 6'h8 == _T_248 ? _GEN_19 : _GEN_1194;
  assign _GEN_1259 = 6'h9 == _T_248 ? _GEN_19 : _GEN_1195;
  assign _GEN_1260 = 6'ha == _T_248 ? _GEN_19 : _GEN_1196;
  assign _GEN_1261 = 6'hb == _T_248 ? _GEN_19 : _GEN_1197;
  assign _GEN_1262 = 6'hc == _T_248 ? _GEN_19 : _GEN_1198;
  assign _GEN_1263 = 6'hd == _T_248 ? _GEN_19 : _GEN_1199;
  assign _GEN_1264 = 6'he == _T_248 ? _GEN_19 : _GEN_1200;
  assign _GEN_1265 = 6'hf == _T_248 ? _GEN_19 : _GEN_1201;
  assign _GEN_1266 = 6'h10 == _T_248 ? _GEN_19 : _GEN_1202;
  assign _GEN_1267 = 6'h11 == _T_248 ? _GEN_19 : _GEN_1203;
  assign _GEN_1268 = 6'h12 == _T_248 ? _GEN_19 : _GEN_1204;
  assign _GEN_1269 = 6'h13 == _T_248 ? _GEN_19 : _GEN_1205;
  assign _GEN_1270 = 6'h14 == _T_248 ? _GEN_19 : _GEN_1206;
  assign _GEN_1271 = 6'h15 == _T_248 ? _GEN_19 : _GEN_1207;
  assign _GEN_1272 = 6'h16 == _T_248 ? _GEN_19 : _GEN_1208;
  assign _GEN_1273 = 6'h17 == _T_248 ? _GEN_19 : _GEN_1209;
  assign _GEN_1274 = 6'h18 == _T_248 ? _GEN_19 : _GEN_1210;
  assign _GEN_1275 = 6'h19 == _T_248 ? _GEN_19 : _GEN_1211;
  assign _GEN_1276 = 6'h1a == _T_248 ? _GEN_19 : _GEN_1212;
  assign _GEN_1277 = 6'h1b == _T_248 ? _GEN_19 : _GEN_1213;
  assign _GEN_1278 = 6'h1c == _T_248 ? _GEN_19 : _GEN_1214;
  assign _GEN_1279 = 6'h1d == _T_248 ? _GEN_19 : _GEN_1215;
  assign _GEN_1280 = 6'h1e == _T_248 ? _GEN_19 : _GEN_1216;
  assign _GEN_1281 = 6'h1f == _T_248 ? _GEN_19 : _GEN_1217;
  assign _GEN_1282 = 6'h20 == _T_248 ? _GEN_19 : _GEN_1218;
  assign _GEN_1283 = 6'h21 == _T_248 ? _GEN_19 : _GEN_1219;
  assign _GEN_1284 = 6'h22 == _T_248 ? _GEN_19 : _GEN_1220;
  assign _GEN_1285 = 6'h23 == _T_248 ? _GEN_19 : _GEN_1221;
  assign _GEN_1286 = 6'h24 == _T_248 ? _GEN_19 : _GEN_1222;
  assign _GEN_1287 = 6'h25 == _T_248 ? _GEN_19 : _GEN_1223;
  assign _GEN_1288 = 6'h26 == _T_248 ? _GEN_19 : _GEN_1224;
  assign _GEN_1289 = 6'h27 == _T_248 ? _GEN_19 : _GEN_1225;
  assign _GEN_1290 = 6'h28 == _T_248 ? _GEN_19 : _GEN_1226;
  assign _GEN_1291 = 6'h29 == _T_248 ? _GEN_19 : _GEN_1227;
  assign _GEN_1292 = 6'h2a == _T_248 ? _GEN_19 : _GEN_1228;
  assign _GEN_1293 = 6'h2b == _T_248 ? _GEN_19 : _GEN_1229;
  assign _GEN_1294 = 6'h2c == _T_248 ? _GEN_19 : _GEN_1230;
  assign _GEN_1295 = 6'h2d == _T_248 ? _GEN_19 : _GEN_1231;
  assign _GEN_1296 = 6'h2e == _T_248 ? _GEN_19 : _GEN_1232;
  assign _GEN_1297 = 6'h2f == _T_248 ? _GEN_19 : _GEN_1233;
  assign _GEN_1298 = 6'h30 == _T_248 ? _GEN_19 : _GEN_1234;
  assign _GEN_1299 = 6'h31 == _T_248 ? _GEN_19 : _GEN_1235;
  assign _GEN_1300 = 6'h32 == _T_248 ? _GEN_19 : _GEN_1236;
  assign _GEN_1301 = 6'h33 == _T_248 ? _GEN_19 : _GEN_1237;
  assign _GEN_1302 = 6'h34 == _T_248 ? _GEN_19 : _GEN_1238;
  assign _GEN_1303 = 6'h35 == _T_248 ? _GEN_19 : _GEN_1239;
  assign _GEN_1304 = 6'h36 == _T_248 ? _GEN_19 : _GEN_1240;
  assign _GEN_1305 = 6'h37 == _T_248 ? _GEN_19 : _GEN_1241;
  assign _GEN_1306 = 6'h38 == _T_248 ? _GEN_19 : _GEN_1242;
  assign _GEN_1307 = 6'h39 == _T_248 ? _GEN_19 : _GEN_1243;
  assign _GEN_1308 = 6'h3a == _T_248 ? _GEN_19 : _GEN_1244;
  assign _GEN_1309 = 6'h3b == _T_248 ? _GEN_19 : _GEN_1245;
  assign _GEN_1310 = 6'h3c == _T_248 ? _GEN_19 : _GEN_1246;
  assign _GEN_1311 = 6'h3d == _T_248 ? _GEN_19 : _GEN_1247;
  assign _GEN_1312 = 6'h3e == _T_248 ? _GEN_19 : _GEN_1248;
  assign _GEN_1313 = 6'h3f == _T_248 ? _GEN_19 : _GEN_1249;
  assign _T_252 = wPos + 6'h14;
  assign _T_253 = _T_252[5:0];
  assign _T_255 = io_fastin[47:44];
  assign _GEN_20 = _T_255;
  assign _GEN_1314 = 6'h0 == _T_253 ? _GEN_20 : _GEN_1250;
  assign _GEN_1315 = 6'h1 == _T_253 ? _GEN_20 : _GEN_1251;
  assign _GEN_1316 = 6'h2 == _T_253 ? _GEN_20 : _GEN_1252;
  assign _GEN_1317 = 6'h3 == _T_253 ? _GEN_20 : _GEN_1253;
  assign _GEN_1318 = 6'h4 == _T_253 ? _GEN_20 : _GEN_1254;
  assign _GEN_1319 = 6'h5 == _T_253 ? _GEN_20 : _GEN_1255;
  assign _GEN_1320 = 6'h6 == _T_253 ? _GEN_20 : _GEN_1256;
  assign _GEN_1321 = 6'h7 == _T_253 ? _GEN_20 : _GEN_1257;
  assign _GEN_1322 = 6'h8 == _T_253 ? _GEN_20 : _GEN_1258;
  assign _GEN_1323 = 6'h9 == _T_253 ? _GEN_20 : _GEN_1259;
  assign _GEN_1324 = 6'ha == _T_253 ? _GEN_20 : _GEN_1260;
  assign _GEN_1325 = 6'hb == _T_253 ? _GEN_20 : _GEN_1261;
  assign _GEN_1326 = 6'hc == _T_253 ? _GEN_20 : _GEN_1262;
  assign _GEN_1327 = 6'hd == _T_253 ? _GEN_20 : _GEN_1263;
  assign _GEN_1328 = 6'he == _T_253 ? _GEN_20 : _GEN_1264;
  assign _GEN_1329 = 6'hf == _T_253 ? _GEN_20 : _GEN_1265;
  assign _GEN_1330 = 6'h10 == _T_253 ? _GEN_20 : _GEN_1266;
  assign _GEN_1331 = 6'h11 == _T_253 ? _GEN_20 : _GEN_1267;
  assign _GEN_1332 = 6'h12 == _T_253 ? _GEN_20 : _GEN_1268;
  assign _GEN_1333 = 6'h13 == _T_253 ? _GEN_20 : _GEN_1269;
  assign _GEN_1334 = 6'h14 == _T_253 ? _GEN_20 : _GEN_1270;
  assign _GEN_1335 = 6'h15 == _T_253 ? _GEN_20 : _GEN_1271;
  assign _GEN_1336 = 6'h16 == _T_253 ? _GEN_20 : _GEN_1272;
  assign _GEN_1337 = 6'h17 == _T_253 ? _GEN_20 : _GEN_1273;
  assign _GEN_1338 = 6'h18 == _T_253 ? _GEN_20 : _GEN_1274;
  assign _GEN_1339 = 6'h19 == _T_253 ? _GEN_20 : _GEN_1275;
  assign _GEN_1340 = 6'h1a == _T_253 ? _GEN_20 : _GEN_1276;
  assign _GEN_1341 = 6'h1b == _T_253 ? _GEN_20 : _GEN_1277;
  assign _GEN_1342 = 6'h1c == _T_253 ? _GEN_20 : _GEN_1278;
  assign _GEN_1343 = 6'h1d == _T_253 ? _GEN_20 : _GEN_1279;
  assign _GEN_1344 = 6'h1e == _T_253 ? _GEN_20 : _GEN_1280;
  assign _GEN_1345 = 6'h1f == _T_253 ? _GEN_20 : _GEN_1281;
  assign _GEN_1346 = 6'h20 == _T_253 ? _GEN_20 : _GEN_1282;
  assign _GEN_1347 = 6'h21 == _T_253 ? _GEN_20 : _GEN_1283;
  assign _GEN_1348 = 6'h22 == _T_253 ? _GEN_20 : _GEN_1284;
  assign _GEN_1349 = 6'h23 == _T_253 ? _GEN_20 : _GEN_1285;
  assign _GEN_1350 = 6'h24 == _T_253 ? _GEN_20 : _GEN_1286;
  assign _GEN_1351 = 6'h25 == _T_253 ? _GEN_20 : _GEN_1287;
  assign _GEN_1352 = 6'h26 == _T_253 ? _GEN_20 : _GEN_1288;
  assign _GEN_1353 = 6'h27 == _T_253 ? _GEN_20 : _GEN_1289;
  assign _GEN_1354 = 6'h28 == _T_253 ? _GEN_20 : _GEN_1290;
  assign _GEN_1355 = 6'h29 == _T_253 ? _GEN_20 : _GEN_1291;
  assign _GEN_1356 = 6'h2a == _T_253 ? _GEN_20 : _GEN_1292;
  assign _GEN_1357 = 6'h2b == _T_253 ? _GEN_20 : _GEN_1293;
  assign _GEN_1358 = 6'h2c == _T_253 ? _GEN_20 : _GEN_1294;
  assign _GEN_1359 = 6'h2d == _T_253 ? _GEN_20 : _GEN_1295;
  assign _GEN_1360 = 6'h2e == _T_253 ? _GEN_20 : _GEN_1296;
  assign _GEN_1361 = 6'h2f == _T_253 ? _GEN_20 : _GEN_1297;
  assign _GEN_1362 = 6'h30 == _T_253 ? _GEN_20 : _GEN_1298;
  assign _GEN_1363 = 6'h31 == _T_253 ? _GEN_20 : _GEN_1299;
  assign _GEN_1364 = 6'h32 == _T_253 ? _GEN_20 : _GEN_1300;
  assign _GEN_1365 = 6'h33 == _T_253 ? _GEN_20 : _GEN_1301;
  assign _GEN_1366 = 6'h34 == _T_253 ? _GEN_20 : _GEN_1302;
  assign _GEN_1367 = 6'h35 == _T_253 ? _GEN_20 : _GEN_1303;
  assign _GEN_1368 = 6'h36 == _T_253 ? _GEN_20 : _GEN_1304;
  assign _GEN_1369 = 6'h37 == _T_253 ? _GEN_20 : _GEN_1305;
  assign _GEN_1370 = 6'h38 == _T_253 ? _GEN_20 : _GEN_1306;
  assign _GEN_1371 = 6'h39 == _T_253 ? _GEN_20 : _GEN_1307;
  assign _GEN_1372 = 6'h3a == _T_253 ? _GEN_20 : _GEN_1308;
  assign _GEN_1373 = 6'h3b == _T_253 ? _GEN_20 : _GEN_1309;
  assign _GEN_1374 = 6'h3c == _T_253 ? _GEN_20 : _GEN_1310;
  assign _GEN_1375 = 6'h3d == _T_253 ? _GEN_20 : _GEN_1311;
  assign _GEN_1376 = 6'h3e == _T_253 ? _GEN_20 : _GEN_1312;
  assign _GEN_1377 = 6'h3f == _T_253 ? _GEN_20 : _GEN_1313;
  assign _T_257 = wPos + 6'h15;
  assign _T_258 = _T_257[5:0];
  assign _T_260 = io_fastin[43:40];
  assign _GEN_21 = _T_260;
  assign _GEN_1378 = 6'h0 == _T_258 ? _GEN_21 : _GEN_1314;
  assign _GEN_1379 = 6'h1 == _T_258 ? _GEN_21 : _GEN_1315;
  assign _GEN_1380 = 6'h2 == _T_258 ? _GEN_21 : _GEN_1316;
  assign _GEN_1381 = 6'h3 == _T_258 ? _GEN_21 : _GEN_1317;
  assign _GEN_1382 = 6'h4 == _T_258 ? _GEN_21 : _GEN_1318;
  assign _GEN_1383 = 6'h5 == _T_258 ? _GEN_21 : _GEN_1319;
  assign _GEN_1384 = 6'h6 == _T_258 ? _GEN_21 : _GEN_1320;
  assign _GEN_1385 = 6'h7 == _T_258 ? _GEN_21 : _GEN_1321;
  assign _GEN_1386 = 6'h8 == _T_258 ? _GEN_21 : _GEN_1322;
  assign _GEN_1387 = 6'h9 == _T_258 ? _GEN_21 : _GEN_1323;
  assign _GEN_1388 = 6'ha == _T_258 ? _GEN_21 : _GEN_1324;
  assign _GEN_1389 = 6'hb == _T_258 ? _GEN_21 : _GEN_1325;
  assign _GEN_1390 = 6'hc == _T_258 ? _GEN_21 : _GEN_1326;
  assign _GEN_1391 = 6'hd == _T_258 ? _GEN_21 : _GEN_1327;
  assign _GEN_1392 = 6'he == _T_258 ? _GEN_21 : _GEN_1328;
  assign _GEN_1393 = 6'hf == _T_258 ? _GEN_21 : _GEN_1329;
  assign _GEN_1394 = 6'h10 == _T_258 ? _GEN_21 : _GEN_1330;
  assign _GEN_1395 = 6'h11 == _T_258 ? _GEN_21 : _GEN_1331;
  assign _GEN_1396 = 6'h12 == _T_258 ? _GEN_21 : _GEN_1332;
  assign _GEN_1397 = 6'h13 == _T_258 ? _GEN_21 : _GEN_1333;
  assign _GEN_1398 = 6'h14 == _T_258 ? _GEN_21 : _GEN_1334;
  assign _GEN_1399 = 6'h15 == _T_258 ? _GEN_21 : _GEN_1335;
  assign _GEN_1400 = 6'h16 == _T_258 ? _GEN_21 : _GEN_1336;
  assign _GEN_1401 = 6'h17 == _T_258 ? _GEN_21 : _GEN_1337;
  assign _GEN_1402 = 6'h18 == _T_258 ? _GEN_21 : _GEN_1338;
  assign _GEN_1403 = 6'h19 == _T_258 ? _GEN_21 : _GEN_1339;
  assign _GEN_1404 = 6'h1a == _T_258 ? _GEN_21 : _GEN_1340;
  assign _GEN_1405 = 6'h1b == _T_258 ? _GEN_21 : _GEN_1341;
  assign _GEN_1406 = 6'h1c == _T_258 ? _GEN_21 : _GEN_1342;
  assign _GEN_1407 = 6'h1d == _T_258 ? _GEN_21 : _GEN_1343;
  assign _GEN_1408 = 6'h1e == _T_258 ? _GEN_21 : _GEN_1344;
  assign _GEN_1409 = 6'h1f == _T_258 ? _GEN_21 : _GEN_1345;
  assign _GEN_1410 = 6'h20 == _T_258 ? _GEN_21 : _GEN_1346;
  assign _GEN_1411 = 6'h21 == _T_258 ? _GEN_21 : _GEN_1347;
  assign _GEN_1412 = 6'h22 == _T_258 ? _GEN_21 : _GEN_1348;
  assign _GEN_1413 = 6'h23 == _T_258 ? _GEN_21 : _GEN_1349;
  assign _GEN_1414 = 6'h24 == _T_258 ? _GEN_21 : _GEN_1350;
  assign _GEN_1415 = 6'h25 == _T_258 ? _GEN_21 : _GEN_1351;
  assign _GEN_1416 = 6'h26 == _T_258 ? _GEN_21 : _GEN_1352;
  assign _GEN_1417 = 6'h27 == _T_258 ? _GEN_21 : _GEN_1353;
  assign _GEN_1418 = 6'h28 == _T_258 ? _GEN_21 : _GEN_1354;
  assign _GEN_1419 = 6'h29 == _T_258 ? _GEN_21 : _GEN_1355;
  assign _GEN_1420 = 6'h2a == _T_258 ? _GEN_21 : _GEN_1356;
  assign _GEN_1421 = 6'h2b == _T_258 ? _GEN_21 : _GEN_1357;
  assign _GEN_1422 = 6'h2c == _T_258 ? _GEN_21 : _GEN_1358;
  assign _GEN_1423 = 6'h2d == _T_258 ? _GEN_21 : _GEN_1359;
  assign _GEN_1424 = 6'h2e == _T_258 ? _GEN_21 : _GEN_1360;
  assign _GEN_1425 = 6'h2f == _T_258 ? _GEN_21 : _GEN_1361;
  assign _GEN_1426 = 6'h30 == _T_258 ? _GEN_21 : _GEN_1362;
  assign _GEN_1427 = 6'h31 == _T_258 ? _GEN_21 : _GEN_1363;
  assign _GEN_1428 = 6'h32 == _T_258 ? _GEN_21 : _GEN_1364;
  assign _GEN_1429 = 6'h33 == _T_258 ? _GEN_21 : _GEN_1365;
  assign _GEN_1430 = 6'h34 == _T_258 ? _GEN_21 : _GEN_1366;
  assign _GEN_1431 = 6'h35 == _T_258 ? _GEN_21 : _GEN_1367;
  assign _GEN_1432 = 6'h36 == _T_258 ? _GEN_21 : _GEN_1368;
  assign _GEN_1433 = 6'h37 == _T_258 ? _GEN_21 : _GEN_1369;
  assign _GEN_1434 = 6'h38 == _T_258 ? _GEN_21 : _GEN_1370;
  assign _GEN_1435 = 6'h39 == _T_258 ? _GEN_21 : _GEN_1371;
  assign _GEN_1436 = 6'h3a == _T_258 ? _GEN_21 : _GEN_1372;
  assign _GEN_1437 = 6'h3b == _T_258 ? _GEN_21 : _GEN_1373;
  assign _GEN_1438 = 6'h3c == _T_258 ? _GEN_21 : _GEN_1374;
  assign _GEN_1439 = 6'h3d == _T_258 ? _GEN_21 : _GEN_1375;
  assign _GEN_1440 = 6'h3e == _T_258 ? _GEN_21 : _GEN_1376;
  assign _GEN_1441 = 6'h3f == _T_258 ? _GEN_21 : _GEN_1377;
  assign _T_262 = wPos + 6'h16;
  assign _T_263 = _T_262[5:0];
  assign _T_265 = io_fastin[39:36];
  assign _GEN_22 = _T_265;
  assign _GEN_1442 = 6'h0 == _T_263 ? _GEN_22 : _GEN_1378;
  assign _GEN_1443 = 6'h1 == _T_263 ? _GEN_22 : _GEN_1379;
  assign _GEN_1444 = 6'h2 == _T_263 ? _GEN_22 : _GEN_1380;
  assign _GEN_1445 = 6'h3 == _T_263 ? _GEN_22 : _GEN_1381;
  assign _GEN_1446 = 6'h4 == _T_263 ? _GEN_22 : _GEN_1382;
  assign _GEN_1447 = 6'h5 == _T_263 ? _GEN_22 : _GEN_1383;
  assign _GEN_1448 = 6'h6 == _T_263 ? _GEN_22 : _GEN_1384;
  assign _GEN_1449 = 6'h7 == _T_263 ? _GEN_22 : _GEN_1385;
  assign _GEN_1450 = 6'h8 == _T_263 ? _GEN_22 : _GEN_1386;
  assign _GEN_1451 = 6'h9 == _T_263 ? _GEN_22 : _GEN_1387;
  assign _GEN_1452 = 6'ha == _T_263 ? _GEN_22 : _GEN_1388;
  assign _GEN_1453 = 6'hb == _T_263 ? _GEN_22 : _GEN_1389;
  assign _GEN_1454 = 6'hc == _T_263 ? _GEN_22 : _GEN_1390;
  assign _GEN_1455 = 6'hd == _T_263 ? _GEN_22 : _GEN_1391;
  assign _GEN_1456 = 6'he == _T_263 ? _GEN_22 : _GEN_1392;
  assign _GEN_1457 = 6'hf == _T_263 ? _GEN_22 : _GEN_1393;
  assign _GEN_1458 = 6'h10 == _T_263 ? _GEN_22 : _GEN_1394;
  assign _GEN_1459 = 6'h11 == _T_263 ? _GEN_22 : _GEN_1395;
  assign _GEN_1460 = 6'h12 == _T_263 ? _GEN_22 : _GEN_1396;
  assign _GEN_1461 = 6'h13 == _T_263 ? _GEN_22 : _GEN_1397;
  assign _GEN_1462 = 6'h14 == _T_263 ? _GEN_22 : _GEN_1398;
  assign _GEN_1463 = 6'h15 == _T_263 ? _GEN_22 : _GEN_1399;
  assign _GEN_1464 = 6'h16 == _T_263 ? _GEN_22 : _GEN_1400;
  assign _GEN_1465 = 6'h17 == _T_263 ? _GEN_22 : _GEN_1401;
  assign _GEN_1466 = 6'h18 == _T_263 ? _GEN_22 : _GEN_1402;
  assign _GEN_1467 = 6'h19 == _T_263 ? _GEN_22 : _GEN_1403;
  assign _GEN_1468 = 6'h1a == _T_263 ? _GEN_22 : _GEN_1404;
  assign _GEN_1469 = 6'h1b == _T_263 ? _GEN_22 : _GEN_1405;
  assign _GEN_1470 = 6'h1c == _T_263 ? _GEN_22 : _GEN_1406;
  assign _GEN_1471 = 6'h1d == _T_263 ? _GEN_22 : _GEN_1407;
  assign _GEN_1472 = 6'h1e == _T_263 ? _GEN_22 : _GEN_1408;
  assign _GEN_1473 = 6'h1f == _T_263 ? _GEN_22 : _GEN_1409;
  assign _GEN_1474 = 6'h20 == _T_263 ? _GEN_22 : _GEN_1410;
  assign _GEN_1475 = 6'h21 == _T_263 ? _GEN_22 : _GEN_1411;
  assign _GEN_1476 = 6'h22 == _T_263 ? _GEN_22 : _GEN_1412;
  assign _GEN_1477 = 6'h23 == _T_263 ? _GEN_22 : _GEN_1413;
  assign _GEN_1478 = 6'h24 == _T_263 ? _GEN_22 : _GEN_1414;
  assign _GEN_1479 = 6'h25 == _T_263 ? _GEN_22 : _GEN_1415;
  assign _GEN_1480 = 6'h26 == _T_263 ? _GEN_22 : _GEN_1416;
  assign _GEN_1481 = 6'h27 == _T_263 ? _GEN_22 : _GEN_1417;
  assign _GEN_1482 = 6'h28 == _T_263 ? _GEN_22 : _GEN_1418;
  assign _GEN_1483 = 6'h29 == _T_263 ? _GEN_22 : _GEN_1419;
  assign _GEN_1484 = 6'h2a == _T_263 ? _GEN_22 : _GEN_1420;
  assign _GEN_1485 = 6'h2b == _T_263 ? _GEN_22 : _GEN_1421;
  assign _GEN_1486 = 6'h2c == _T_263 ? _GEN_22 : _GEN_1422;
  assign _GEN_1487 = 6'h2d == _T_263 ? _GEN_22 : _GEN_1423;
  assign _GEN_1488 = 6'h2e == _T_263 ? _GEN_22 : _GEN_1424;
  assign _GEN_1489 = 6'h2f == _T_263 ? _GEN_22 : _GEN_1425;
  assign _GEN_1490 = 6'h30 == _T_263 ? _GEN_22 : _GEN_1426;
  assign _GEN_1491 = 6'h31 == _T_263 ? _GEN_22 : _GEN_1427;
  assign _GEN_1492 = 6'h32 == _T_263 ? _GEN_22 : _GEN_1428;
  assign _GEN_1493 = 6'h33 == _T_263 ? _GEN_22 : _GEN_1429;
  assign _GEN_1494 = 6'h34 == _T_263 ? _GEN_22 : _GEN_1430;
  assign _GEN_1495 = 6'h35 == _T_263 ? _GEN_22 : _GEN_1431;
  assign _GEN_1496 = 6'h36 == _T_263 ? _GEN_22 : _GEN_1432;
  assign _GEN_1497 = 6'h37 == _T_263 ? _GEN_22 : _GEN_1433;
  assign _GEN_1498 = 6'h38 == _T_263 ? _GEN_22 : _GEN_1434;
  assign _GEN_1499 = 6'h39 == _T_263 ? _GEN_22 : _GEN_1435;
  assign _GEN_1500 = 6'h3a == _T_263 ? _GEN_22 : _GEN_1436;
  assign _GEN_1501 = 6'h3b == _T_263 ? _GEN_22 : _GEN_1437;
  assign _GEN_1502 = 6'h3c == _T_263 ? _GEN_22 : _GEN_1438;
  assign _GEN_1503 = 6'h3d == _T_263 ? _GEN_22 : _GEN_1439;
  assign _GEN_1504 = 6'h3e == _T_263 ? _GEN_22 : _GEN_1440;
  assign _GEN_1505 = 6'h3f == _T_263 ? _GEN_22 : _GEN_1441;
  assign _T_267 = wPos + 6'h17;
  assign _T_268 = _T_267[5:0];
  assign _T_270 = io_fastin[35:32];
  assign _GEN_23 = _T_270;
  assign _GEN_1506 = 6'h0 == _T_268 ? _GEN_23 : _GEN_1442;
  assign _GEN_1507 = 6'h1 == _T_268 ? _GEN_23 : _GEN_1443;
  assign _GEN_1508 = 6'h2 == _T_268 ? _GEN_23 : _GEN_1444;
  assign _GEN_1509 = 6'h3 == _T_268 ? _GEN_23 : _GEN_1445;
  assign _GEN_1510 = 6'h4 == _T_268 ? _GEN_23 : _GEN_1446;
  assign _GEN_1511 = 6'h5 == _T_268 ? _GEN_23 : _GEN_1447;
  assign _GEN_1512 = 6'h6 == _T_268 ? _GEN_23 : _GEN_1448;
  assign _GEN_1513 = 6'h7 == _T_268 ? _GEN_23 : _GEN_1449;
  assign _GEN_1514 = 6'h8 == _T_268 ? _GEN_23 : _GEN_1450;
  assign _GEN_1515 = 6'h9 == _T_268 ? _GEN_23 : _GEN_1451;
  assign _GEN_1516 = 6'ha == _T_268 ? _GEN_23 : _GEN_1452;
  assign _GEN_1517 = 6'hb == _T_268 ? _GEN_23 : _GEN_1453;
  assign _GEN_1518 = 6'hc == _T_268 ? _GEN_23 : _GEN_1454;
  assign _GEN_1519 = 6'hd == _T_268 ? _GEN_23 : _GEN_1455;
  assign _GEN_1520 = 6'he == _T_268 ? _GEN_23 : _GEN_1456;
  assign _GEN_1521 = 6'hf == _T_268 ? _GEN_23 : _GEN_1457;
  assign _GEN_1522 = 6'h10 == _T_268 ? _GEN_23 : _GEN_1458;
  assign _GEN_1523 = 6'h11 == _T_268 ? _GEN_23 : _GEN_1459;
  assign _GEN_1524 = 6'h12 == _T_268 ? _GEN_23 : _GEN_1460;
  assign _GEN_1525 = 6'h13 == _T_268 ? _GEN_23 : _GEN_1461;
  assign _GEN_1526 = 6'h14 == _T_268 ? _GEN_23 : _GEN_1462;
  assign _GEN_1527 = 6'h15 == _T_268 ? _GEN_23 : _GEN_1463;
  assign _GEN_1528 = 6'h16 == _T_268 ? _GEN_23 : _GEN_1464;
  assign _GEN_1529 = 6'h17 == _T_268 ? _GEN_23 : _GEN_1465;
  assign _GEN_1530 = 6'h18 == _T_268 ? _GEN_23 : _GEN_1466;
  assign _GEN_1531 = 6'h19 == _T_268 ? _GEN_23 : _GEN_1467;
  assign _GEN_1532 = 6'h1a == _T_268 ? _GEN_23 : _GEN_1468;
  assign _GEN_1533 = 6'h1b == _T_268 ? _GEN_23 : _GEN_1469;
  assign _GEN_1534 = 6'h1c == _T_268 ? _GEN_23 : _GEN_1470;
  assign _GEN_1535 = 6'h1d == _T_268 ? _GEN_23 : _GEN_1471;
  assign _GEN_1536 = 6'h1e == _T_268 ? _GEN_23 : _GEN_1472;
  assign _GEN_1537 = 6'h1f == _T_268 ? _GEN_23 : _GEN_1473;
  assign _GEN_1538 = 6'h20 == _T_268 ? _GEN_23 : _GEN_1474;
  assign _GEN_1539 = 6'h21 == _T_268 ? _GEN_23 : _GEN_1475;
  assign _GEN_1540 = 6'h22 == _T_268 ? _GEN_23 : _GEN_1476;
  assign _GEN_1541 = 6'h23 == _T_268 ? _GEN_23 : _GEN_1477;
  assign _GEN_1542 = 6'h24 == _T_268 ? _GEN_23 : _GEN_1478;
  assign _GEN_1543 = 6'h25 == _T_268 ? _GEN_23 : _GEN_1479;
  assign _GEN_1544 = 6'h26 == _T_268 ? _GEN_23 : _GEN_1480;
  assign _GEN_1545 = 6'h27 == _T_268 ? _GEN_23 : _GEN_1481;
  assign _GEN_1546 = 6'h28 == _T_268 ? _GEN_23 : _GEN_1482;
  assign _GEN_1547 = 6'h29 == _T_268 ? _GEN_23 : _GEN_1483;
  assign _GEN_1548 = 6'h2a == _T_268 ? _GEN_23 : _GEN_1484;
  assign _GEN_1549 = 6'h2b == _T_268 ? _GEN_23 : _GEN_1485;
  assign _GEN_1550 = 6'h2c == _T_268 ? _GEN_23 : _GEN_1486;
  assign _GEN_1551 = 6'h2d == _T_268 ? _GEN_23 : _GEN_1487;
  assign _GEN_1552 = 6'h2e == _T_268 ? _GEN_23 : _GEN_1488;
  assign _GEN_1553 = 6'h2f == _T_268 ? _GEN_23 : _GEN_1489;
  assign _GEN_1554 = 6'h30 == _T_268 ? _GEN_23 : _GEN_1490;
  assign _GEN_1555 = 6'h31 == _T_268 ? _GEN_23 : _GEN_1491;
  assign _GEN_1556 = 6'h32 == _T_268 ? _GEN_23 : _GEN_1492;
  assign _GEN_1557 = 6'h33 == _T_268 ? _GEN_23 : _GEN_1493;
  assign _GEN_1558 = 6'h34 == _T_268 ? _GEN_23 : _GEN_1494;
  assign _GEN_1559 = 6'h35 == _T_268 ? _GEN_23 : _GEN_1495;
  assign _GEN_1560 = 6'h36 == _T_268 ? _GEN_23 : _GEN_1496;
  assign _GEN_1561 = 6'h37 == _T_268 ? _GEN_23 : _GEN_1497;
  assign _GEN_1562 = 6'h38 == _T_268 ? _GEN_23 : _GEN_1498;
  assign _GEN_1563 = 6'h39 == _T_268 ? _GEN_23 : _GEN_1499;
  assign _GEN_1564 = 6'h3a == _T_268 ? _GEN_23 : _GEN_1500;
  assign _GEN_1565 = 6'h3b == _T_268 ? _GEN_23 : _GEN_1501;
  assign _GEN_1566 = 6'h3c == _T_268 ? _GEN_23 : _GEN_1502;
  assign _GEN_1567 = 6'h3d == _T_268 ? _GEN_23 : _GEN_1503;
  assign _GEN_1568 = 6'h3e == _T_268 ? _GEN_23 : _GEN_1504;
  assign _GEN_1569 = 6'h3f == _T_268 ? _GEN_23 : _GEN_1505;
  assign _T_272 = wPos + 6'h18;
  assign _T_273 = _T_272[5:0];
  assign _T_275 = io_fastin[31:28];
  assign _GEN_24 = _T_275;
  assign _GEN_1570 = 6'h0 == _T_273 ? _GEN_24 : _GEN_1506;
  assign _GEN_1571 = 6'h1 == _T_273 ? _GEN_24 : _GEN_1507;
  assign _GEN_1572 = 6'h2 == _T_273 ? _GEN_24 : _GEN_1508;
  assign _GEN_1573 = 6'h3 == _T_273 ? _GEN_24 : _GEN_1509;
  assign _GEN_1574 = 6'h4 == _T_273 ? _GEN_24 : _GEN_1510;
  assign _GEN_1575 = 6'h5 == _T_273 ? _GEN_24 : _GEN_1511;
  assign _GEN_1576 = 6'h6 == _T_273 ? _GEN_24 : _GEN_1512;
  assign _GEN_1577 = 6'h7 == _T_273 ? _GEN_24 : _GEN_1513;
  assign _GEN_1578 = 6'h8 == _T_273 ? _GEN_24 : _GEN_1514;
  assign _GEN_1579 = 6'h9 == _T_273 ? _GEN_24 : _GEN_1515;
  assign _GEN_1580 = 6'ha == _T_273 ? _GEN_24 : _GEN_1516;
  assign _GEN_1581 = 6'hb == _T_273 ? _GEN_24 : _GEN_1517;
  assign _GEN_1582 = 6'hc == _T_273 ? _GEN_24 : _GEN_1518;
  assign _GEN_1583 = 6'hd == _T_273 ? _GEN_24 : _GEN_1519;
  assign _GEN_1584 = 6'he == _T_273 ? _GEN_24 : _GEN_1520;
  assign _GEN_1585 = 6'hf == _T_273 ? _GEN_24 : _GEN_1521;
  assign _GEN_1586 = 6'h10 == _T_273 ? _GEN_24 : _GEN_1522;
  assign _GEN_1587 = 6'h11 == _T_273 ? _GEN_24 : _GEN_1523;
  assign _GEN_1588 = 6'h12 == _T_273 ? _GEN_24 : _GEN_1524;
  assign _GEN_1589 = 6'h13 == _T_273 ? _GEN_24 : _GEN_1525;
  assign _GEN_1590 = 6'h14 == _T_273 ? _GEN_24 : _GEN_1526;
  assign _GEN_1591 = 6'h15 == _T_273 ? _GEN_24 : _GEN_1527;
  assign _GEN_1592 = 6'h16 == _T_273 ? _GEN_24 : _GEN_1528;
  assign _GEN_1593 = 6'h17 == _T_273 ? _GEN_24 : _GEN_1529;
  assign _GEN_1594 = 6'h18 == _T_273 ? _GEN_24 : _GEN_1530;
  assign _GEN_1595 = 6'h19 == _T_273 ? _GEN_24 : _GEN_1531;
  assign _GEN_1596 = 6'h1a == _T_273 ? _GEN_24 : _GEN_1532;
  assign _GEN_1597 = 6'h1b == _T_273 ? _GEN_24 : _GEN_1533;
  assign _GEN_1598 = 6'h1c == _T_273 ? _GEN_24 : _GEN_1534;
  assign _GEN_1599 = 6'h1d == _T_273 ? _GEN_24 : _GEN_1535;
  assign _GEN_1600 = 6'h1e == _T_273 ? _GEN_24 : _GEN_1536;
  assign _GEN_1601 = 6'h1f == _T_273 ? _GEN_24 : _GEN_1537;
  assign _GEN_1602 = 6'h20 == _T_273 ? _GEN_24 : _GEN_1538;
  assign _GEN_1603 = 6'h21 == _T_273 ? _GEN_24 : _GEN_1539;
  assign _GEN_1604 = 6'h22 == _T_273 ? _GEN_24 : _GEN_1540;
  assign _GEN_1605 = 6'h23 == _T_273 ? _GEN_24 : _GEN_1541;
  assign _GEN_1606 = 6'h24 == _T_273 ? _GEN_24 : _GEN_1542;
  assign _GEN_1607 = 6'h25 == _T_273 ? _GEN_24 : _GEN_1543;
  assign _GEN_1608 = 6'h26 == _T_273 ? _GEN_24 : _GEN_1544;
  assign _GEN_1609 = 6'h27 == _T_273 ? _GEN_24 : _GEN_1545;
  assign _GEN_1610 = 6'h28 == _T_273 ? _GEN_24 : _GEN_1546;
  assign _GEN_1611 = 6'h29 == _T_273 ? _GEN_24 : _GEN_1547;
  assign _GEN_1612 = 6'h2a == _T_273 ? _GEN_24 : _GEN_1548;
  assign _GEN_1613 = 6'h2b == _T_273 ? _GEN_24 : _GEN_1549;
  assign _GEN_1614 = 6'h2c == _T_273 ? _GEN_24 : _GEN_1550;
  assign _GEN_1615 = 6'h2d == _T_273 ? _GEN_24 : _GEN_1551;
  assign _GEN_1616 = 6'h2e == _T_273 ? _GEN_24 : _GEN_1552;
  assign _GEN_1617 = 6'h2f == _T_273 ? _GEN_24 : _GEN_1553;
  assign _GEN_1618 = 6'h30 == _T_273 ? _GEN_24 : _GEN_1554;
  assign _GEN_1619 = 6'h31 == _T_273 ? _GEN_24 : _GEN_1555;
  assign _GEN_1620 = 6'h32 == _T_273 ? _GEN_24 : _GEN_1556;
  assign _GEN_1621 = 6'h33 == _T_273 ? _GEN_24 : _GEN_1557;
  assign _GEN_1622 = 6'h34 == _T_273 ? _GEN_24 : _GEN_1558;
  assign _GEN_1623 = 6'h35 == _T_273 ? _GEN_24 : _GEN_1559;
  assign _GEN_1624 = 6'h36 == _T_273 ? _GEN_24 : _GEN_1560;
  assign _GEN_1625 = 6'h37 == _T_273 ? _GEN_24 : _GEN_1561;
  assign _GEN_1626 = 6'h38 == _T_273 ? _GEN_24 : _GEN_1562;
  assign _GEN_1627 = 6'h39 == _T_273 ? _GEN_24 : _GEN_1563;
  assign _GEN_1628 = 6'h3a == _T_273 ? _GEN_24 : _GEN_1564;
  assign _GEN_1629 = 6'h3b == _T_273 ? _GEN_24 : _GEN_1565;
  assign _GEN_1630 = 6'h3c == _T_273 ? _GEN_24 : _GEN_1566;
  assign _GEN_1631 = 6'h3d == _T_273 ? _GEN_24 : _GEN_1567;
  assign _GEN_1632 = 6'h3e == _T_273 ? _GEN_24 : _GEN_1568;
  assign _GEN_1633 = 6'h3f == _T_273 ? _GEN_24 : _GEN_1569;
  assign _T_277 = wPos + 6'h19;
  assign _T_278 = _T_277[5:0];
  assign _T_280 = io_fastin[27:24];
  assign _GEN_25 = _T_280;
  assign _GEN_1634 = 6'h0 == _T_278 ? _GEN_25 : _GEN_1570;
  assign _GEN_1635 = 6'h1 == _T_278 ? _GEN_25 : _GEN_1571;
  assign _GEN_1636 = 6'h2 == _T_278 ? _GEN_25 : _GEN_1572;
  assign _GEN_1637 = 6'h3 == _T_278 ? _GEN_25 : _GEN_1573;
  assign _GEN_1638 = 6'h4 == _T_278 ? _GEN_25 : _GEN_1574;
  assign _GEN_1639 = 6'h5 == _T_278 ? _GEN_25 : _GEN_1575;
  assign _GEN_1640 = 6'h6 == _T_278 ? _GEN_25 : _GEN_1576;
  assign _GEN_1641 = 6'h7 == _T_278 ? _GEN_25 : _GEN_1577;
  assign _GEN_1642 = 6'h8 == _T_278 ? _GEN_25 : _GEN_1578;
  assign _GEN_1643 = 6'h9 == _T_278 ? _GEN_25 : _GEN_1579;
  assign _GEN_1644 = 6'ha == _T_278 ? _GEN_25 : _GEN_1580;
  assign _GEN_1645 = 6'hb == _T_278 ? _GEN_25 : _GEN_1581;
  assign _GEN_1646 = 6'hc == _T_278 ? _GEN_25 : _GEN_1582;
  assign _GEN_1647 = 6'hd == _T_278 ? _GEN_25 : _GEN_1583;
  assign _GEN_1648 = 6'he == _T_278 ? _GEN_25 : _GEN_1584;
  assign _GEN_1649 = 6'hf == _T_278 ? _GEN_25 : _GEN_1585;
  assign _GEN_1650 = 6'h10 == _T_278 ? _GEN_25 : _GEN_1586;
  assign _GEN_1651 = 6'h11 == _T_278 ? _GEN_25 : _GEN_1587;
  assign _GEN_1652 = 6'h12 == _T_278 ? _GEN_25 : _GEN_1588;
  assign _GEN_1653 = 6'h13 == _T_278 ? _GEN_25 : _GEN_1589;
  assign _GEN_1654 = 6'h14 == _T_278 ? _GEN_25 : _GEN_1590;
  assign _GEN_1655 = 6'h15 == _T_278 ? _GEN_25 : _GEN_1591;
  assign _GEN_1656 = 6'h16 == _T_278 ? _GEN_25 : _GEN_1592;
  assign _GEN_1657 = 6'h17 == _T_278 ? _GEN_25 : _GEN_1593;
  assign _GEN_1658 = 6'h18 == _T_278 ? _GEN_25 : _GEN_1594;
  assign _GEN_1659 = 6'h19 == _T_278 ? _GEN_25 : _GEN_1595;
  assign _GEN_1660 = 6'h1a == _T_278 ? _GEN_25 : _GEN_1596;
  assign _GEN_1661 = 6'h1b == _T_278 ? _GEN_25 : _GEN_1597;
  assign _GEN_1662 = 6'h1c == _T_278 ? _GEN_25 : _GEN_1598;
  assign _GEN_1663 = 6'h1d == _T_278 ? _GEN_25 : _GEN_1599;
  assign _GEN_1664 = 6'h1e == _T_278 ? _GEN_25 : _GEN_1600;
  assign _GEN_1665 = 6'h1f == _T_278 ? _GEN_25 : _GEN_1601;
  assign _GEN_1666 = 6'h20 == _T_278 ? _GEN_25 : _GEN_1602;
  assign _GEN_1667 = 6'h21 == _T_278 ? _GEN_25 : _GEN_1603;
  assign _GEN_1668 = 6'h22 == _T_278 ? _GEN_25 : _GEN_1604;
  assign _GEN_1669 = 6'h23 == _T_278 ? _GEN_25 : _GEN_1605;
  assign _GEN_1670 = 6'h24 == _T_278 ? _GEN_25 : _GEN_1606;
  assign _GEN_1671 = 6'h25 == _T_278 ? _GEN_25 : _GEN_1607;
  assign _GEN_1672 = 6'h26 == _T_278 ? _GEN_25 : _GEN_1608;
  assign _GEN_1673 = 6'h27 == _T_278 ? _GEN_25 : _GEN_1609;
  assign _GEN_1674 = 6'h28 == _T_278 ? _GEN_25 : _GEN_1610;
  assign _GEN_1675 = 6'h29 == _T_278 ? _GEN_25 : _GEN_1611;
  assign _GEN_1676 = 6'h2a == _T_278 ? _GEN_25 : _GEN_1612;
  assign _GEN_1677 = 6'h2b == _T_278 ? _GEN_25 : _GEN_1613;
  assign _GEN_1678 = 6'h2c == _T_278 ? _GEN_25 : _GEN_1614;
  assign _GEN_1679 = 6'h2d == _T_278 ? _GEN_25 : _GEN_1615;
  assign _GEN_1680 = 6'h2e == _T_278 ? _GEN_25 : _GEN_1616;
  assign _GEN_1681 = 6'h2f == _T_278 ? _GEN_25 : _GEN_1617;
  assign _GEN_1682 = 6'h30 == _T_278 ? _GEN_25 : _GEN_1618;
  assign _GEN_1683 = 6'h31 == _T_278 ? _GEN_25 : _GEN_1619;
  assign _GEN_1684 = 6'h32 == _T_278 ? _GEN_25 : _GEN_1620;
  assign _GEN_1685 = 6'h33 == _T_278 ? _GEN_25 : _GEN_1621;
  assign _GEN_1686 = 6'h34 == _T_278 ? _GEN_25 : _GEN_1622;
  assign _GEN_1687 = 6'h35 == _T_278 ? _GEN_25 : _GEN_1623;
  assign _GEN_1688 = 6'h36 == _T_278 ? _GEN_25 : _GEN_1624;
  assign _GEN_1689 = 6'h37 == _T_278 ? _GEN_25 : _GEN_1625;
  assign _GEN_1690 = 6'h38 == _T_278 ? _GEN_25 : _GEN_1626;
  assign _GEN_1691 = 6'h39 == _T_278 ? _GEN_25 : _GEN_1627;
  assign _GEN_1692 = 6'h3a == _T_278 ? _GEN_25 : _GEN_1628;
  assign _GEN_1693 = 6'h3b == _T_278 ? _GEN_25 : _GEN_1629;
  assign _GEN_1694 = 6'h3c == _T_278 ? _GEN_25 : _GEN_1630;
  assign _GEN_1695 = 6'h3d == _T_278 ? _GEN_25 : _GEN_1631;
  assign _GEN_1696 = 6'h3e == _T_278 ? _GEN_25 : _GEN_1632;
  assign _GEN_1697 = 6'h3f == _T_278 ? _GEN_25 : _GEN_1633;
  assign _T_282 = wPos + 6'h1a;
  assign _T_283 = _T_282[5:0];
  assign _T_285 = io_fastin[23:20];
  assign _GEN_26 = _T_285;
  assign _GEN_1698 = 6'h0 == _T_283 ? _GEN_26 : _GEN_1634;
  assign _GEN_1699 = 6'h1 == _T_283 ? _GEN_26 : _GEN_1635;
  assign _GEN_1700 = 6'h2 == _T_283 ? _GEN_26 : _GEN_1636;
  assign _GEN_1701 = 6'h3 == _T_283 ? _GEN_26 : _GEN_1637;
  assign _GEN_1702 = 6'h4 == _T_283 ? _GEN_26 : _GEN_1638;
  assign _GEN_1703 = 6'h5 == _T_283 ? _GEN_26 : _GEN_1639;
  assign _GEN_1704 = 6'h6 == _T_283 ? _GEN_26 : _GEN_1640;
  assign _GEN_1705 = 6'h7 == _T_283 ? _GEN_26 : _GEN_1641;
  assign _GEN_1706 = 6'h8 == _T_283 ? _GEN_26 : _GEN_1642;
  assign _GEN_1707 = 6'h9 == _T_283 ? _GEN_26 : _GEN_1643;
  assign _GEN_1708 = 6'ha == _T_283 ? _GEN_26 : _GEN_1644;
  assign _GEN_1709 = 6'hb == _T_283 ? _GEN_26 : _GEN_1645;
  assign _GEN_1710 = 6'hc == _T_283 ? _GEN_26 : _GEN_1646;
  assign _GEN_1711 = 6'hd == _T_283 ? _GEN_26 : _GEN_1647;
  assign _GEN_1712 = 6'he == _T_283 ? _GEN_26 : _GEN_1648;
  assign _GEN_1713 = 6'hf == _T_283 ? _GEN_26 : _GEN_1649;
  assign _GEN_1714 = 6'h10 == _T_283 ? _GEN_26 : _GEN_1650;
  assign _GEN_1715 = 6'h11 == _T_283 ? _GEN_26 : _GEN_1651;
  assign _GEN_1716 = 6'h12 == _T_283 ? _GEN_26 : _GEN_1652;
  assign _GEN_1717 = 6'h13 == _T_283 ? _GEN_26 : _GEN_1653;
  assign _GEN_1718 = 6'h14 == _T_283 ? _GEN_26 : _GEN_1654;
  assign _GEN_1719 = 6'h15 == _T_283 ? _GEN_26 : _GEN_1655;
  assign _GEN_1720 = 6'h16 == _T_283 ? _GEN_26 : _GEN_1656;
  assign _GEN_1721 = 6'h17 == _T_283 ? _GEN_26 : _GEN_1657;
  assign _GEN_1722 = 6'h18 == _T_283 ? _GEN_26 : _GEN_1658;
  assign _GEN_1723 = 6'h19 == _T_283 ? _GEN_26 : _GEN_1659;
  assign _GEN_1724 = 6'h1a == _T_283 ? _GEN_26 : _GEN_1660;
  assign _GEN_1725 = 6'h1b == _T_283 ? _GEN_26 : _GEN_1661;
  assign _GEN_1726 = 6'h1c == _T_283 ? _GEN_26 : _GEN_1662;
  assign _GEN_1727 = 6'h1d == _T_283 ? _GEN_26 : _GEN_1663;
  assign _GEN_1728 = 6'h1e == _T_283 ? _GEN_26 : _GEN_1664;
  assign _GEN_1729 = 6'h1f == _T_283 ? _GEN_26 : _GEN_1665;
  assign _GEN_1730 = 6'h20 == _T_283 ? _GEN_26 : _GEN_1666;
  assign _GEN_1731 = 6'h21 == _T_283 ? _GEN_26 : _GEN_1667;
  assign _GEN_1732 = 6'h22 == _T_283 ? _GEN_26 : _GEN_1668;
  assign _GEN_1733 = 6'h23 == _T_283 ? _GEN_26 : _GEN_1669;
  assign _GEN_1734 = 6'h24 == _T_283 ? _GEN_26 : _GEN_1670;
  assign _GEN_1735 = 6'h25 == _T_283 ? _GEN_26 : _GEN_1671;
  assign _GEN_1736 = 6'h26 == _T_283 ? _GEN_26 : _GEN_1672;
  assign _GEN_1737 = 6'h27 == _T_283 ? _GEN_26 : _GEN_1673;
  assign _GEN_1738 = 6'h28 == _T_283 ? _GEN_26 : _GEN_1674;
  assign _GEN_1739 = 6'h29 == _T_283 ? _GEN_26 : _GEN_1675;
  assign _GEN_1740 = 6'h2a == _T_283 ? _GEN_26 : _GEN_1676;
  assign _GEN_1741 = 6'h2b == _T_283 ? _GEN_26 : _GEN_1677;
  assign _GEN_1742 = 6'h2c == _T_283 ? _GEN_26 : _GEN_1678;
  assign _GEN_1743 = 6'h2d == _T_283 ? _GEN_26 : _GEN_1679;
  assign _GEN_1744 = 6'h2e == _T_283 ? _GEN_26 : _GEN_1680;
  assign _GEN_1745 = 6'h2f == _T_283 ? _GEN_26 : _GEN_1681;
  assign _GEN_1746 = 6'h30 == _T_283 ? _GEN_26 : _GEN_1682;
  assign _GEN_1747 = 6'h31 == _T_283 ? _GEN_26 : _GEN_1683;
  assign _GEN_1748 = 6'h32 == _T_283 ? _GEN_26 : _GEN_1684;
  assign _GEN_1749 = 6'h33 == _T_283 ? _GEN_26 : _GEN_1685;
  assign _GEN_1750 = 6'h34 == _T_283 ? _GEN_26 : _GEN_1686;
  assign _GEN_1751 = 6'h35 == _T_283 ? _GEN_26 : _GEN_1687;
  assign _GEN_1752 = 6'h36 == _T_283 ? _GEN_26 : _GEN_1688;
  assign _GEN_1753 = 6'h37 == _T_283 ? _GEN_26 : _GEN_1689;
  assign _GEN_1754 = 6'h38 == _T_283 ? _GEN_26 : _GEN_1690;
  assign _GEN_1755 = 6'h39 == _T_283 ? _GEN_26 : _GEN_1691;
  assign _GEN_1756 = 6'h3a == _T_283 ? _GEN_26 : _GEN_1692;
  assign _GEN_1757 = 6'h3b == _T_283 ? _GEN_26 : _GEN_1693;
  assign _GEN_1758 = 6'h3c == _T_283 ? _GEN_26 : _GEN_1694;
  assign _GEN_1759 = 6'h3d == _T_283 ? _GEN_26 : _GEN_1695;
  assign _GEN_1760 = 6'h3e == _T_283 ? _GEN_26 : _GEN_1696;
  assign _GEN_1761 = 6'h3f == _T_283 ? _GEN_26 : _GEN_1697;
  assign _T_287 = wPos + 6'h1b;
  assign _T_288 = _T_287[5:0];
  assign _T_290 = io_fastin[19:16];
  assign _GEN_27 = _T_290;
  assign _GEN_1762 = 6'h0 == _T_288 ? _GEN_27 : _GEN_1698;
  assign _GEN_1763 = 6'h1 == _T_288 ? _GEN_27 : _GEN_1699;
  assign _GEN_1764 = 6'h2 == _T_288 ? _GEN_27 : _GEN_1700;
  assign _GEN_1765 = 6'h3 == _T_288 ? _GEN_27 : _GEN_1701;
  assign _GEN_1766 = 6'h4 == _T_288 ? _GEN_27 : _GEN_1702;
  assign _GEN_1767 = 6'h5 == _T_288 ? _GEN_27 : _GEN_1703;
  assign _GEN_1768 = 6'h6 == _T_288 ? _GEN_27 : _GEN_1704;
  assign _GEN_1769 = 6'h7 == _T_288 ? _GEN_27 : _GEN_1705;
  assign _GEN_1770 = 6'h8 == _T_288 ? _GEN_27 : _GEN_1706;
  assign _GEN_1771 = 6'h9 == _T_288 ? _GEN_27 : _GEN_1707;
  assign _GEN_1772 = 6'ha == _T_288 ? _GEN_27 : _GEN_1708;
  assign _GEN_1773 = 6'hb == _T_288 ? _GEN_27 : _GEN_1709;
  assign _GEN_1774 = 6'hc == _T_288 ? _GEN_27 : _GEN_1710;
  assign _GEN_1775 = 6'hd == _T_288 ? _GEN_27 : _GEN_1711;
  assign _GEN_1776 = 6'he == _T_288 ? _GEN_27 : _GEN_1712;
  assign _GEN_1777 = 6'hf == _T_288 ? _GEN_27 : _GEN_1713;
  assign _GEN_1778 = 6'h10 == _T_288 ? _GEN_27 : _GEN_1714;
  assign _GEN_1779 = 6'h11 == _T_288 ? _GEN_27 : _GEN_1715;
  assign _GEN_1780 = 6'h12 == _T_288 ? _GEN_27 : _GEN_1716;
  assign _GEN_1781 = 6'h13 == _T_288 ? _GEN_27 : _GEN_1717;
  assign _GEN_1782 = 6'h14 == _T_288 ? _GEN_27 : _GEN_1718;
  assign _GEN_1783 = 6'h15 == _T_288 ? _GEN_27 : _GEN_1719;
  assign _GEN_1784 = 6'h16 == _T_288 ? _GEN_27 : _GEN_1720;
  assign _GEN_1785 = 6'h17 == _T_288 ? _GEN_27 : _GEN_1721;
  assign _GEN_1786 = 6'h18 == _T_288 ? _GEN_27 : _GEN_1722;
  assign _GEN_1787 = 6'h19 == _T_288 ? _GEN_27 : _GEN_1723;
  assign _GEN_1788 = 6'h1a == _T_288 ? _GEN_27 : _GEN_1724;
  assign _GEN_1789 = 6'h1b == _T_288 ? _GEN_27 : _GEN_1725;
  assign _GEN_1790 = 6'h1c == _T_288 ? _GEN_27 : _GEN_1726;
  assign _GEN_1791 = 6'h1d == _T_288 ? _GEN_27 : _GEN_1727;
  assign _GEN_1792 = 6'h1e == _T_288 ? _GEN_27 : _GEN_1728;
  assign _GEN_1793 = 6'h1f == _T_288 ? _GEN_27 : _GEN_1729;
  assign _GEN_1794 = 6'h20 == _T_288 ? _GEN_27 : _GEN_1730;
  assign _GEN_1795 = 6'h21 == _T_288 ? _GEN_27 : _GEN_1731;
  assign _GEN_1796 = 6'h22 == _T_288 ? _GEN_27 : _GEN_1732;
  assign _GEN_1797 = 6'h23 == _T_288 ? _GEN_27 : _GEN_1733;
  assign _GEN_1798 = 6'h24 == _T_288 ? _GEN_27 : _GEN_1734;
  assign _GEN_1799 = 6'h25 == _T_288 ? _GEN_27 : _GEN_1735;
  assign _GEN_1800 = 6'h26 == _T_288 ? _GEN_27 : _GEN_1736;
  assign _GEN_1801 = 6'h27 == _T_288 ? _GEN_27 : _GEN_1737;
  assign _GEN_1802 = 6'h28 == _T_288 ? _GEN_27 : _GEN_1738;
  assign _GEN_1803 = 6'h29 == _T_288 ? _GEN_27 : _GEN_1739;
  assign _GEN_1804 = 6'h2a == _T_288 ? _GEN_27 : _GEN_1740;
  assign _GEN_1805 = 6'h2b == _T_288 ? _GEN_27 : _GEN_1741;
  assign _GEN_1806 = 6'h2c == _T_288 ? _GEN_27 : _GEN_1742;
  assign _GEN_1807 = 6'h2d == _T_288 ? _GEN_27 : _GEN_1743;
  assign _GEN_1808 = 6'h2e == _T_288 ? _GEN_27 : _GEN_1744;
  assign _GEN_1809 = 6'h2f == _T_288 ? _GEN_27 : _GEN_1745;
  assign _GEN_1810 = 6'h30 == _T_288 ? _GEN_27 : _GEN_1746;
  assign _GEN_1811 = 6'h31 == _T_288 ? _GEN_27 : _GEN_1747;
  assign _GEN_1812 = 6'h32 == _T_288 ? _GEN_27 : _GEN_1748;
  assign _GEN_1813 = 6'h33 == _T_288 ? _GEN_27 : _GEN_1749;
  assign _GEN_1814 = 6'h34 == _T_288 ? _GEN_27 : _GEN_1750;
  assign _GEN_1815 = 6'h35 == _T_288 ? _GEN_27 : _GEN_1751;
  assign _GEN_1816 = 6'h36 == _T_288 ? _GEN_27 : _GEN_1752;
  assign _GEN_1817 = 6'h37 == _T_288 ? _GEN_27 : _GEN_1753;
  assign _GEN_1818 = 6'h38 == _T_288 ? _GEN_27 : _GEN_1754;
  assign _GEN_1819 = 6'h39 == _T_288 ? _GEN_27 : _GEN_1755;
  assign _GEN_1820 = 6'h3a == _T_288 ? _GEN_27 : _GEN_1756;
  assign _GEN_1821 = 6'h3b == _T_288 ? _GEN_27 : _GEN_1757;
  assign _GEN_1822 = 6'h3c == _T_288 ? _GEN_27 : _GEN_1758;
  assign _GEN_1823 = 6'h3d == _T_288 ? _GEN_27 : _GEN_1759;
  assign _GEN_1824 = 6'h3e == _T_288 ? _GEN_27 : _GEN_1760;
  assign _GEN_1825 = 6'h3f == _T_288 ? _GEN_27 : _GEN_1761;
  assign _T_292 = wPos + 6'h1c;
  assign _T_293 = _T_292[5:0];
  assign _T_295 = io_fastin[15:12];
  assign _GEN_28 = _T_295;
  assign _GEN_1826 = 6'h0 == _T_293 ? _GEN_28 : _GEN_1762;
  assign _GEN_1827 = 6'h1 == _T_293 ? _GEN_28 : _GEN_1763;
  assign _GEN_1828 = 6'h2 == _T_293 ? _GEN_28 : _GEN_1764;
  assign _GEN_1829 = 6'h3 == _T_293 ? _GEN_28 : _GEN_1765;
  assign _GEN_1830 = 6'h4 == _T_293 ? _GEN_28 : _GEN_1766;
  assign _GEN_1831 = 6'h5 == _T_293 ? _GEN_28 : _GEN_1767;
  assign _GEN_1832 = 6'h6 == _T_293 ? _GEN_28 : _GEN_1768;
  assign _GEN_1833 = 6'h7 == _T_293 ? _GEN_28 : _GEN_1769;
  assign _GEN_1834 = 6'h8 == _T_293 ? _GEN_28 : _GEN_1770;
  assign _GEN_1835 = 6'h9 == _T_293 ? _GEN_28 : _GEN_1771;
  assign _GEN_1836 = 6'ha == _T_293 ? _GEN_28 : _GEN_1772;
  assign _GEN_1837 = 6'hb == _T_293 ? _GEN_28 : _GEN_1773;
  assign _GEN_1838 = 6'hc == _T_293 ? _GEN_28 : _GEN_1774;
  assign _GEN_1839 = 6'hd == _T_293 ? _GEN_28 : _GEN_1775;
  assign _GEN_1840 = 6'he == _T_293 ? _GEN_28 : _GEN_1776;
  assign _GEN_1841 = 6'hf == _T_293 ? _GEN_28 : _GEN_1777;
  assign _GEN_1842 = 6'h10 == _T_293 ? _GEN_28 : _GEN_1778;
  assign _GEN_1843 = 6'h11 == _T_293 ? _GEN_28 : _GEN_1779;
  assign _GEN_1844 = 6'h12 == _T_293 ? _GEN_28 : _GEN_1780;
  assign _GEN_1845 = 6'h13 == _T_293 ? _GEN_28 : _GEN_1781;
  assign _GEN_1846 = 6'h14 == _T_293 ? _GEN_28 : _GEN_1782;
  assign _GEN_1847 = 6'h15 == _T_293 ? _GEN_28 : _GEN_1783;
  assign _GEN_1848 = 6'h16 == _T_293 ? _GEN_28 : _GEN_1784;
  assign _GEN_1849 = 6'h17 == _T_293 ? _GEN_28 : _GEN_1785;
  assign _GEN_1850 = 6'h18 == _T_293 ? _GEN_28 : _GEN_1786;
  assign _GEN_1851 = 6'h19 == _T_293 ? _GEN_28 : _GEN_1787;
  assign _GEN_1852 = 6'h1a == _T_293 ? _GEN_28 : _GEN_1788;
  assign _GEN_1853 = 6'h1b == _T_293 ? _GEN_28 : _GEN_1789;
  assign _GEN_1854 = 6'h1c == _T_293 ? _GEN_28 : _GEN_1790;
  assign _GEN_1855 = 6'h1d == _T_293 ? _GEN_28 : _GEN_1791;
  assign _GEN_1856 = 6'h1e == _T_293 ? _GEN_28 : _GEN_1792;
  assign _GEN_1857 = 6'h1f == _T_293 ? _GEN_28 : _GEN_1793;
  assign _GEN_1858 = 6'h20 == _T_293 ? _GEN_28 : _GEN_1794;
  assign _GEN_1859 = 6'h21 == _T_293 ? _GEN_28 : _GEN_1795;
  assign _GEN_1860 = 6'h22 == _T_293 ? _GEN_28 : _GEN_1796;
  assign _GEN_1861 = 6'h23 == _T_293 ? _GEN_28 : _GEN_1797;
  assign _GEN_1862 = 6'h24 == _T_293 ? _GEN_28 : _GEN_1798;
  assign _GEN_1863 = 6'h25 == _T_293 ? _GEN_28 : _GEN_1799;
  assign _GEN_1864 = 6'h26 == _T_293 ? _GEN_28 : _GEN_1800;
  assign _GEN_1865 = 6'h27 == _T_293 ? _GEN_28 : _GEN_1801;
  assign _GEN_1866 = 6'h28 == _T_293 ? _GEN_28 : _GEN_1802;
  assign _GEN_1867 = 6'h29 == _T_293 ? _GEN_28 : _GEN_1803;
  assign _GEN_1868 = 6'h2a == _T_293 ? _GEN_28 : _GEN_1804;
  assign _GEN_1869 = 6'h2b == _T_293 ? _GEN_28 : _GEN_1805;
  assign _GEN_1870 = 6'h2c == _T_293 ? _GEN_28 : _GEN_1806;
  assign _GEN_1871 = 6'h2d == _T_293 ? _GEN_28 : _GEN_1807;
  assign _GEN_1872 = 6'h2e == _T_293 ? _GEN_28 : _GEN_1808;
  assign _GEN_1873 = 6'h2f == _T_293 ? _GEN_28 : _GEN_1809;
  assign _GEN_1874 = 6'h30 == _T_293 ? _GEN_28 : _GEN_1810;
  assign _GEN_1875 = 6'h31 == _T_293 ? _GEN_28 : _GEN_1811;
  assign _GEN_1876 = 6'h32 == _T_293 ? _GEN_28 : _GEN_1812;
  assign _GEN_1877 = 6'h33 == _T_293 ? _GEN_28 : _GEN_1813;
  assign _GEN_1878 = 6'h34 == _T_293 ? _GEN_28 : _GEN_1814;
  assign _GEN_1879 = 6'h35 == _T_293 ? _GEN_28 : _GEN_1815;
  assign _GEN_1880 = 6'h36 == _T_293 ? _GEN_28 : _GEN_1816;
  assign _GEN_1881 = 6'h37 == _T_293 ? _GEN_28 : _GEN_1817;
  assign _GEN_1882 = 6'h38 == _T_293 ? _GEN_28 : _GEN_1818;
  assign _GEN_1883 = 6'h39 == _T_293 ? _GEN_28 : _GEN_1819;
  assign _GEN_1884 = 6'h3a == _T_293 ? _GEN_28 : _GEN_1820;
  assign _GEN_1885 = 6'h3b == _T_293 ? _GEN_28 : _GEN_1821;
  assign _GEN_1886 = 6'h3c == _T_293 ? _GEN_28 : _GEN_1822;
  assign _GEN_1887 = 6'h3d == _T_293 ? _GEN_28 : _GEN_1823;
  assign _GEN_1888 = 6'h3e == _T_293 ? _GEN_28 : _GEN_1824;
  assign _GEN_1889 = 6'h3f == _T_293 ? _GEN_28 : _GEN_1825;
  assign _T_297 = wPos + 6'h1d;
  assign _T_298 = _T_297[5:0];
  assign _T_300 = io_fastin[11:8];
  assign _GEN_29 = _T_300;
  assign _GEN_1890 = 6'h0 == _T_298 ? _GEN_29 : _GEN_1826;
  assign _GEN_1891 = 6'h1 == _T_298 ? _GEN_29 : _GEN_1827;
  assign _GEN_1892 = 6'h2 == _T_298 ? _GEN_29 : _GEN_1828;
  assign _GEN_1893 = 6'h3 == _T_298 ? _GEN_29 : _GEN_1829;
  assign _GEN_1894 = 6'h4 == _T_298 ? _GEN_29 : _GEN_1830;
  assign _GEN_1895 = 6'h5 == _T_298 ? _GEN_29 : _GEN_1831;
  assign _GEN_1896 = 6'h6 == _T_298 ? _GEN_29 : _GEN_1832;
  assign _GEN_1897 = 6'h7 == _T_298 ? _GEN_29 : _GEN_1833;
  assign _GEN_1898 = 6'h8 == _T_298 ? _GEN_29 : _GEN_1834;
  assign _GEN_1899 = 6'h9 == _T_298 ? _GEN_29 : _GEN_1835;
  assign _GEN_1900 = 6'ha == _T_298 ? _GEN_29 : _GEN_1836;
  assign _GEN_1901 = 6'hb == _T_298 ? _GEN_29 : _GEN_1837;
  assign _GEN_1902 = 6'hc == _T_298 ? _GEN_29 : _GEN_1838;
  assign _GEN_1903 = 6'hd == _T_298 ? _GEN_29 : _GEN_1839;
  assign _GEN_1904 = 6'he == _T_298 ? _GEN_29 : _GEN_1840;
  assign _GEN_1905 = 6'hf == _T_298 ? _GEN_29 : _GEN_1841;
  assign _GEN_1906 = 6'h10 == _T_298 ? _GEN_29 : _GEN_1842;
  assign _GEN_1907 = 6'h11 == _T_298 ? _GEN_29 : _GEN_1843;
  assign _GEN_1908 = 6'h12 == _T_298 ? _GEN_29 : _GEN_1844;
  assign _GEN_1909 = 6'h13 == _T_298 ? _GEN_29 : _GEN_1845;
  assign _GEN_1910 = 6'h14 == _T_298 ? _GEN_29 : _GEN_1846;
  assign _GEN_1911 = 6'h15 == _T_298 ? _GEN_29 : _GEN_1847;
  assign _GEN_1912 = 6'h16 == _T_298 ? _GEN_29 : _GEN_1848;
  assign _GEN_1913 = 6'h17 == _T_298 ? _GEN_29 : _GEN_1849;
  assign _GEN_1914 = 6'h18 == _T_298 ? _GEN_29 : _GEN_1850;
  assign _GEN_1915 = 6'h19 == _T_298 ? _GEN_29 : _GEN_1851;
  assign _GEN_1916 = 6'h1a == _T_298 ? _GEN_29 : _GEN_1852;
  assign _GEN_1917 = 6'h1b == _T_298 ? _GEN_29 : _GEN_1853;
  assign _GEN_1918 = 6'h1c == _T_298 ? _GEN_29 : _GEN_1854;
  assign _GEN_1919 = 6'h1d == _T_298 ? _GEN_29 : _GEN_1855;
  assign _GEN_1920 = 6'h1e == _T_298 ? _GEN_29 : _GEN_1856;
  assign _GEN_1921 = 6'h1f == _T_298 ? _GEN_29 : _GEN_1857;
  assign _GEN_1922 = 6'h20 == _T_298 ? _GEN_29 : _GEN_1858;
  assign _GEN_1923 = 6'h21 == _T_298 ? _GEN_29 : _GEN_1859;
  assign _GEN_1924 = 6'h22 == _T_298 ? _GEN_29 : _GEN_1860;
  assign _GEN_1925 = 6'h23 == _T_298 ? _GEN_29 : _GEN_1861;
  assign _GEN_1926 = 6'h24 == _T_298 ? _GEN_29 : _GEN_1862;
  assign _GEN_1927 = 6'h25 == _T_298 ? _GEN_29 : _GEN_1863;
  assign _GEN_1928 = 6'h26 == _T_298 ? _GEN_29 : _GEN_1864;
  assign _GEN_1929 = 6'h27 == _T_298 ? _GEN_29 : _GEN_1865;
  assign _GEN_1930 = 6'h28 == _T_298 ? _GEN_29 : _GEN_1866;
  assign _GEN_1931 = 6'h29 == _T_298 ? _GEN_29 : _GEN_1867;
  assign _GEN_1932 = 6'h2a == _T_298 ? _GEN_29 : _GEN_1868;
  assign _GEN_1933 = 6'h2b == _T_298 ? _GEN_29 : _GEN_1869;
  assign _GEN_1934 = 6'h2c == _T_298 ? _GEN_29 : _GEN_1870;
  assign _GEN_1935 = 6'h2d == _T_298 ? _GEN_29 : _GEN_1871;
  assign _GEN_1936 = 6'h2e == _T_298 ? _GEN_29 : _GEN_1872;
  assign _GEN_1937 = 6'h2f == _T_298 ? _GEN_29 : _GEN_1873;
  assign _GEN_1938 = 6'h30 == _T_298 ? _GEN_29 : _GEN_1874;
  assign _GEN_1939 = 6'h31 == _T_298 ? _GEN_29 : _GEN_1875;
  assign _GEN_1940 = 6'h32 == _T_298 ? _GEN_29 : _GEN_1876;
  assign _GEN_1941 = 6'h33 == _T_298 ? _GEN_29 : _GEN_1877;
  assign _GEN_1942 = 6'h34 == _T_298 ? _GEN_29 : _GEN_1878;
  assign _GEN_1943 = 6'h35 == _T_298 ? _GEN_29 : _GEN_1879;
  assign _GEN_1944 = 6'h36 == _T_298 ? _GEN_29 : _GEN_1880;
  assign _GEN_1945 = 6'h37 == _T_298 ? _GEN_29 : _GEN_1881;
  assign _GEN_1946 = 6'h38 == _T_298 ? _GEN_29 : _GEN_1882;
  assign _GEN_1947 = 6'h39 == _T_298 ? _GEN_29 : _GEN_1883;
  assign _GEN_1948 = 6'h3a == _T_298 ? _GEN_29 : _GEN_1884;
  assign _GEN_1949 = 6'h3b == _T_298 ? _GEN_29 : _GEN_1885;
  assign _GEN_1950 = 6'h3c == _T_298 ? _GEN_29 : _GEN_1886;
  assign _GEN_1951 = 6'h3d == _T_298 ? _GEN_29 : _GEN_1887;
  assign _GEN_1952 = 6'h3e == _T_298 ? _GEN_29 : _GEN_1888;
  assign _GEN_1953 = 6'h3f == _T_298 ? _GEN_29 : _GEN_1889;
  assign _T_302 = wPos + 6'h1e;
  assign _T_303 = _T_302[5:0];
  assign _T_305 = io_fastin[7:4];
  assign _GEN_30 = _T_305;
  assign _GEN_1954 = 6'h0 == _T_303 ? _GEN_30 : _GEN_1890;
  assign _GEN_1955 = 6'h1 == _T_303 ? _GEN_30 : _GEN_1891;
  assign _GEN_1956 = 6'h2 == _T_303 ? _GEN_30 : _GEN_1892;
  assign _GEN_1957 = 6'h3 == _T_303 ? _GEN_30 : _GEN_1893;
  assign _GEN_1958 = 6'h4 == _T_303 ? _GEN_30 : _GEN_1894;
  assign _GEN_1959 = 6'h5 == _T_303 ? _GEN_30 : _GEN_1895;
  assign _GEN_1960 = 6'h6 == _T_303 ? _GEN_30 : _GEN_1896;
  assign _GEN_1961 = 6'h7 == _T_303 ? _GEN_30 : _GEN_1897;
  assign _GEN_1962 = 6'h8 == _T_303 ? _GEN_30 : _GEN_1898;
  assign _GEN_1963 = 6'h9 == _T_303 ? _GEN_30 : _GEN_1899;
  assign _GEN_1964 = 6'ha == _T_303 ? _GEN_30 : _GEN_1900;
  assign _GEN_1965 = 6'hb == _T_303 ? _GEN_30 : _GEN_1901;
  assign _GEN_1966 = 6'hc == _T_303 ? _GEN_30 : _GEN_1902;
  assign _GEN_1967 = 6'hd == _T_303 ? _GEN_30 : _GEN_1903;
  assign _GEN_1968 = 6'he == _T_303 ? _GEN_30 : _GEN_1904;
  assign _GEN_1969 = 6'hf == _T_303 ? _GEN_30 : _GEN_1905;
  assign _GEN_1970 = 6'h10 == _T_303 ? _GEN_30 : _GEN_1906;
  assign _GEN_1971 = 6'h11 == _T_303 ? _GEN_30 : _GEN_1907;
  assign _GEN_1972 = 6'h12 == _T_303 ? _GEN_30 : _GEN_1908;
  assign _GEN_1973 = 6'h13 == _T_303 ? _GEN_30 : _GEN_1909;
  assign _GEN_1974 = 6'h14 == _T_303 ? _GEN_30 : _GEN_1910;
  assign _GEN_1975 = 6'h15 == _T_303 ? _GEN_30 : _GEN_1911;
  assign _GEN_1976 = 6'h16 == _T_303 ? _GEN_30 : _GEN_1912;
  assign _GEN_1977 = 6'h17 == _T_303 ? _GEN_30 : _GEN_1913;
  assign _GEN_1978 = 6'h18 == _T_303 ? _GEN_30 : _GEN_1914;
  assign _GEN_1979 = 6'h19 == _T_303 ? _GEN_30 : _GEN_1915;
  assign _GEN_1980 = 6'h1a == _T_303 ? _GEN_30 : _GEN_1916;
  assign _GEN_1981 = 6'h1b == _T_303 ? _GEN_30 : _GEN_1917;
  assign _GEN_1982 = 6'h1c == _T_303 ? _GEN_30 : _GEN_1918;
  assign _GEN_1983 = 6'h1d == _T_303 ? _GEN_30 : _GEN_1919;
  assign _GEN_1984 = 6'h1e == _T_303 ? _GEN_30 : _GEN_1920;
  assign _GEN_1985 = 6'h1f == _T_303 ? _GEN_30 : _GEN_1921;
  assign _GEN_1986 = 6'h20 == _T_303 ? _GEN_30 : _GEN_1922;
  assign _GEN_1987 = 6'h21 == _T_303 ? _GEN_30 : _GEN_1923;
  assign _GEN_1988 = 6'h22 == _T_303 ? _GEN_30 : _GEN_1924;
  assign _GEN_1989 = 6'h23 == _T_303 ? _GEN_30 : _GEN_1925;
  assign _GEN_1990 = 6'h24 == _T_303 ? _GEN_30 : _GEN_1926;
  assign _GEN_1991 = 6'h25 == _T_303 ? _GEN_30 : _GEN_1927;
  assign _GEN_1992 = 6'h26 == _T_303 ? _GEN_30 : _GEN_1928;
  assign _GEN_1993 = 6'h27 == _T_303 ? _GEN_30 : _GEN_1929;
  assign _GEN_1994 = 6'h28 == _T_303 ? _GEN_30 : _GEN_1930;
  assign _GEN_1995 = 6'h29 == _T_303 ? _GEN_30 : _GEN_1931;
  assign _GEN_1996 = 6'h2a == _T_303 ? _GEN_30 : _GEN_1932;
  assign _GEN_1997 = 6'h2b == _T_303 ? _GEN_30 : _GEN_1933;
  assign _GEN_1998 = 6'h2c == _T_303 ? _GEN_30 : _GEN_1934;
  assign _GEN_1999 = 6'h2d == _T_303 ? _GEN_30 : _GEN_1935;
  assign _GEN_2000 = 6'h2e == _T_303 ? _GEN_30 : _GEN_1936;
  assign _GEN_2001 = 6'h2f == _T_303 ? _GEN_30 : _GEN_1937;
  assign _GEN_2002 = 6'h30 == _T_303 ? _GEN_30 : _GEN_1938;
  assign _GEN_2003 = 6'h31 == _T_303 ? _GEN_30 : _GEN_1939;
  assign _GEN_2004 = 6'h32 == _T_303 ? _GEN_30 : _GEN_1940;
  assign _GEN_2005 = 6'h33 == _T_303 ? _GEN_30 : _GEN_1941;
  assign _GEN_2006 = 6'h34 == _T_303 ? _GEN_30 : _GEN_1942;
  assign _GEN_2007 = 6'h35 == _T_303 ? _GEN_30 : _GEN_1943;
  assign _GEN_2008 = 6'h36 == _T_303 ? _GEN_30 : _GEN_1944;
  assign _GEN_2009 = 6'h37 == _T_303 ? _GEN_30 : _GEN_1945;
  assign _GEN_2010 = 6'h38 == _T_303 ? _GEN_30 : _GEN_1946;
  assign _GEN_2011 = 6'h39 == _T_303 ? _GEN_30 : _GEN_1947;
  assign _GEN_2012 = 6'h3a == _T_303 ? _GEN_30 : _GEN_1948;
  assign _GEN_2013 = 6'h3b == _T_303 ? _GEN_30 : _GEN_1949;
  assign _GEN_2014 = 6'h3c == _T_303 ? _GEN_30 : _GEN_1950;
  assign _GEN_2015 = 6'h3d == _T_303 ? _GEN_30 : _GEN_1951;
  assign _GEN_2016 = 6'h3e == _T_303 ? _GEN_30 : _GEN_1952;
  assign _GEN_2017 = 6'h3f == _T_303 ? _GEN_30 : _GEN_1953;
  assign _T_307 = wPos + 6'h1f;
  assign _T_308 = _T_307[5:0];
  assign _T_310 = io_fastin[3:0];
  assign _GEN_31 = _T_310;
  assign _GEN_2018 = 6'h0 == _T_308 ? _GEN_31 : _GEN_1954;
  assign _GEN_2019 = 6'h1 == _T_308 ? _GEN_31 : _GEN_1955;
  assign _GEN_2020 = 6'h2 == _T_308 ? _GEN_31 : _GEN_1956;
  assign _GEN_2021 = 6'h3 == _T_308 ? _GEN_31 : _GEN_1957;
  assign _GEN_2022 = 6'h4 == _T_308 ? _GEN_31 : _GEN_1958;
  assign _GEN_2023 = 6'h5 == _T_308 ? _GEN_31 : _GEN_1959;
  assign _GEN_2024 = 6'h6 == _T_308 ? _GEN_31 : _GEN_1960;
  assign _GEN_2025 = 6'h7 == _T_308 ? _GEN_31 : _GEN_1961;
  assign _GEN_2026 = 6'h8 == _T_308 ? _GEN_31 : _GEN_1962;
  assign _GEN_2027 = 6'h9 == _T_308 ? _GEN_31 : _GEN_1963;
  assign _GEN_2028 = 6'ha == _T_308 ? _GEN_31 : _GEN_1964;
  assign _GEN_2029 = 6'hb == _T_308 ? _GEN_31 : _GEN_1965;
  assign _GEN_2030 = 6'hc == _T_308 ? _GEN_31 : _GEN_1966;
  assign _GEN_2031 = 6'hd == _T_308 ? _GEN_31 : _GEN_1967;
  assign _GEN_2032 = 6'he == _T_308 ? _GEN_31 : _GEN_1968;
  assign _GEN_2033 = 6'hf == _T_308 ? _GEN_31 : _GEN_1969;
  assign _GEN_2034 = 6'h10 == _T_308 ? _GEN_31 : _GEN_1970;
  assign _GEN_2035 = 6'h11 == _T_308 ? _GEN_31 : _GEN_1971;
  assign _GEN_2036 = 6'h12 == _T_308 ? _GEN_31 : _GEN_1972;
  assign _GEN_2037 = 6'h13 == _T_308 ? _GEN_31 : _GEN_1973;
  assign _GEN_2038 = 6'h14 == _T_308 ? _GEN_31 : _GEN_1974;
  assign _GEN_2039 = 6'h15 == _T_308 ? _GEN_31 : _GEN_1975;
  assign _GEN_2040 = 6'h16 == _T_308 ? _GEN_31 : _GEN_1976;
  assign _GEN_2041 = 6'h17 == _T_308 ? _GEN_31 : _GEN_1977;
  assign _GEN_2042 = 6'h18 == _T_308 ? _GEN_31 : _GEN_1978;
  assign _GEN_2043 = 6'h19 == _T_308 ? _GEN_31 : _GEN_1979;
  assign _GEN_2044 = 6'h1a == _T_308 ? _GEN_31 : _GEN_1980;
  assign _GEN_2045 = 6'h1b == _T_308 ? _GEN_31 : _GEN_1981;
  assign _GEN_2046 = 6'h1c == _T_308 ? _GEN_31 : _GEN_1982;
  assign _GEN_2047 = 6'h1d == _T_308 ? _GEN_31 : _GEN_1983;
  assign _GEN_2048 = 6'h1e == _T_308 ? _GEN_31 : _GEN_1984;
  assign _GEN_2049 = 6'h1f == _T_308 ? _GEN_31 : _GEN_1985;
  assign _GEN_2050 = 6'h20 == _T_308 ? _GEN_31 : _GEN_1986;
  assign _GEN_2051 = 6'h21 == _T_308 ? _GEN_31 : _GEN_1987;
  assign _GEN_2052 = 6'h22 == _T_308 ? _GEN_31 : _GEN_1988;
  assign _GEN_2053 = 6'h23 == _T_308 ? _GEN_31 : _GEN_1989;
  assign _GEN_2054 = 6'h24 == _T_308 ? _GEN_31 : _GEN_1990;
  assign _GEN_2055 = 6'h25 == _T_308 ? _GEN_31 : _GEN_1991;
  assign _GEN_2056 = 6'h26 == _T_308 ? _GEN_31 : _GEN_1992;
  assign _GEN_2057 = 6'h27 == _T_308 ? _GEN_31 : _GEN_1993;
  assign _GEN_2058 = 6'h28 == _T_308 ? _GEN_31 : _GEN_1994;
  assign _GEN_2059 = 6'h29 == _T_308 ? _GEN_31 : _GEN_1995;
  assign _GEN_2060 = 6'h2a == _T_308 ? _GEN_31 : _GEN_1996;
  assign _GEN_2061 = 6'h2b == _T_308 ? _GEN_31 : _GEN_1997;
  assign _GEN_2062 = 6'h2c == _T_308 ? _GEN_31 : _GEN_1998;
  assign _GEN_2063 = 6'h2d == _T_308 ? _GEN_31 : _GEN_1999;
  assign _GEN_2064 = 6'h2e == _T_308 ? _GEN_31 : _GEN_2000;
  assign _GEN_2065 = 6'h2f == _T_308 ? _GEN_31 : _GEN_2001;
  assign _GEN_2066 = 6'h30 == _T_308 ? _GEN_31 : _GEN_2002;
  assign _GEN_2067 = 6'h31 == _T_308 ? _GEN_31 : _GEN_2003;
  assign _GEN_2068 = 6'h32 == _T_308 ? _GEN_31 : _GEN_2004;
  assign _GEN_2069 = 6'h33 == _T_308 ? _GEN_31 : _GEN_2005;
  assign _GEN_2070 = 6'h34 == _T_308 ? _GEN_31 : _GEN_2006;
  assign _GEN_2071 = 6'h35 == _T_308 ? _GEN_31 : _GEN_2007;
  assign _GEN_2072 = 6'h36 == _T_308 ? _GEN_31 : _GEN_2008;
  assign _GEN_2073 = 6'h37 == _T_308 ? _GEN_31 : _GEN_2009;
  assign _GEN_2074 = 6'h38 == _T_308 ? _GEN_31 : _GEN_2010;
  assign _GEN_2075 = 6'h39 == _T_308 ? _GEN_31 : _GEN_2011;
  assign _GEN_2076 = 6'h3a == _T_308 ? _GEN_31 : _GEN_2012;
  assign _GEN_2077 = 6'h3b == _T_308 ? _GEN_31 : _GEN_2013;
  assign _GEN_2078 = 6'h3c == _T_308 ? _GEN_31 : _GEN_2014;
  assign _GEN_2079 = 6'h3d == _T_308 ? _GEN_31 : _GEN_2015;
  assign _GEN_2080 = 6'h3e == _T_308 ? _GEN_31 : _GEN_2016;
  assign _GEN_2081 = 6'h3f == _T_308 ? _GEN_31 : _GEN_2017;
  assign _T_312 = wPos + 6'h20;
  assign _T_313 = _T_312[5:0];
  assign _GEN_2082 = _T_150 ? _GEN_2018 : mem_0;
  assign _GEN_2083 = _T_150 ? _GEN_2019 : mem_1;
  assign _GEN_2084 = _T_150 ? _GEN_2020 : mem_2;
  assign _GEN_2085 = _T_150 ? _GEN_2021 : mem_3;
  assign _GEN_2086 = _T_150 ? _GEN_2022 : mem_4;
  assign _GEN_2087 = _T_150 ? _GEN_2023 : mem_5;
  assign _GEN_2088 = _T_150 ? _GEN_2024 : mem_6;
  assign _GEN_2089 = _T_150 ? _GEN_2025 : mem_7;
  assign _GEN_2090 = _T_150 ? _GEN_2026 : mem_8;
  assign _GEN_2091 = _T_150 ? _GEN_2027 : mem_9;
  assign _GEN_2092 = _T_150 ? _GEN_2028 : mem_10;
  assign _GEN_2093 = _T_150 ? _GEN_2029 : mem_11;
  assign _GEN_2094 = _T_150 ? _GEN_2030 : mem_12;
  assign _GEN_2095 = _T_150 ? _GEN_2031 : mem_13;
  assign _GEN_2096 = _T_150 ? _GEN_2032 : mem_14;
  assign _GEN_2097 = _T_150 ? _GEN_2033 : mem_15;
  assign _GEN_2098 = _T_150 ? _GEN_2034 : mem_16;
  assign _GEN_2099 = _T_150 ? _GEN_2035 : mem_17;
  assign _GEN_2100 = _T_150 ? _GEN_2036 : mem_18;
  assign _GEN_2101 = _T_150 ? _GEN_2037 : mem_19;
  assign _GEN_2102 = _T_150 ? _GEN_2038 : mem_20;
  assign _GEN_2103 = _T_150 ? _GEN_2039 : mem_21;
  assign _GEN_2104 = _T_150 ? _GEN_2040 : mem_22;
  assign _GEN_2105 = _T_150 ? _GEN_2041 : mem_23;
  assign _GEN_2106 = _T_150 ? _GEN_2042 : mem_24;
  assign _GEN_2107 = _T_150 ? _GEN_2043 : mem_25;
  assign _GEN_2108 = _T_150 ? _GEN_2044 : mem_26;
  assign _GEN_2109 = _T_150 ? _GEN_2045 : mem_27;
  assign _GEN_2110 = _T_150 ? _GEN_2046 : mem_28;
  assign _GEN_2111 = _T_150 ? _GEN_2047 : mem_29;
  assign _GEN_2112 = _T_150 ? _GEN_2048 : mem_30;
  assign _GEN_2113 = _T_150 ? _GEN_2049 : mem_31;
  assign _GEN_2114 = _T_150 ? _GEN_2050 : mem_32;
  assign _GEN_2115 = _T_150 ? _GEN_2051 : mem_33;
  assign _GEN_2116 = _T_150 ? _GEN_2052 : mem_34;
  assign _GEN_2117 = _T_150 ? _GEN_2053 : mem_35;
  assign _GEN_2118 = _T_150 ? _GEN_2054 : mem_36;
  assign _GEN_2119 = _T_150 ? _GEN_2055 : mem_37;
  assign _GEN_2120 = _T_150 ? _GEN_2056 : mem_38;
  assign _GEN_2121 = _T_150 ? _GEN_2057 : mem_39;
  assign _GEN_2122 = _T_150 ? _GEN_2058 : mem_40;
  assign _GEN_2123 = _T_150 ? _GEN_2059 : mem_41;
  assign _GEN_2124 = _T_150 ? _GEN_2060 : mem_42;
  assign _GEN_2125 = _T_150 ? _GEN_2061 : mem_43;
  assign _GEN_2126 = _T_150 ? _GEN_2062 : mem_44;
  assign _GEN_2127 = _T_150 ? _GEN_2063 : mem_45;
  assign _GEN_2128 = _T_150 ? _GEN_2064 : mem_46;
  assign _GEN_2129 = _T_150 ? _GEN_2065 : mem_47;
  assign _GEN_2130 = _T_150 ? _GEN_2066 : mem_48;
  assign _GEN_2131 = _T_150 ? _GEN_2067 : mem_49;
  assign _GEN_2132 = _T_150 ? _GEN_2068 : mem_50;
  assign _GEN_2133 = _T_150 ? _GEN_2069 : mem_51;
  assign _GEN_2134 = _T_150 ? _GEN_2070 : mem_52;
  assign _GEN_2135 = _T_150 ? _GEN_2071 : mem_53;
  assign _GEN_2136 = _T_150 ? _GEN_2072 : mem_54;
  assign _GEN_2137 = _T_150 ? _GEN_2073 : mem_55;
  assign _GEN_2138 = _T_150 ? _GEN_2074 : mem_56;
  assign _GEN_2139 = _T_150 ? _GEN_2075 : mem_57;
  assign _GEN_2140 = _T_150 ? _GEN_2076 : mem_58;
  assign _GEN_2141 = _T_150 ? _GEN_2077 : mem_59;
  assign _GEN_2142 = _T_150 ? _GEN_2078 : mem_60;
  assign _GEN_2143 = _T_150 ? _GEN_2079 : mem_61;
  assign _GEN_2144 = _T_150 ? _GEN_2080 : mem_62;
  assign _GEN_2145 = _T_150 ? _GEN_2081 : mem_63;
  assign _GEN_2146 = _T_150 ? _T_313 : wPos;
  assign _T_315 = _T_150 == 1'h0;
  assign _GEN_32 = io_in;
  assign _GEN_2147 = 6'h0 == wPos ? _GEN_32 : _GEN_2082;
  assign _GEN_2148 = 6'h1 == wPos ? _GEN_32 : _GEN_2083;
  assign _GEN_2149 = 6'h2 == wPos ? _GEN_32 : _GEN_2084;
  assign _GEN_2150 = 6'h3 == wPos ? _GEN_32 : _GEN_2085;
  assign _GEN_2151 = 6'h4 == wPos ? _GEN_32 : _GEN_2086;
  assign _GEN_2152 = 6'h5 == wPos ? _GEN_32 : _GEN_2087;
  assign _GEN_2153 = 6'h6 == wPos ? _GEN_32 : _GEN_2088;
  assign _GEN_2154 = 6'h7 == wPos ? _GEN_32 : _GEN_2089;
  assign _GEN_2155 = 6'h8 == wPos ? _GEN_32 : _GEN_2090;
  assign _GEN_2156 = 6'h9 == wPos ? _GEN_32 : _GEN_2091;
  assign _GEN_2157 = 6'ha == wPos ? _GEN_32 : _GEN_2092;
  assign _GEN_2158 = 6'hb == wPos ? _GEN_32 : _GEN_2093;
  assign _GEN_2159 = 6'hc == wPos ? _GEN_32 : _GEN_2094;
  assign _GEN_2160 = 6'hd == wPos ? _GEN_32 : _GEN_2095;
  assign _GEN_2161 = 6'he == wPos ? _GEN_32 : _GEN_2096;
  assign _GEN_2162 = 6'hf == wPos ? _GEN_32 : _GEN_2097;
  assign _GEN_2163 = 6'h10 == wPos ? _GEN_32 : _GEN_2098;
  assign _GEN_2164 = 6'h11 == wPos ? _GEN_32 : _GEN_2099;
  assign _GEN_2165 = 6'h12 == wPos ? _GEN_32 : _GEN_2100;
  assign _GEN_2166 = 6'h13 == wPos ? _GEN_32 : _GEN_2101;
  assign _GEN_2167 = 6'h14 == wPos ? _GEN_32 : _GEN_2102;
  assign _GEN_2168 = 6'h15 == wPos ? _GEN_32 : _GEN_2103;
  assign _GEN_2169 = 6'h16 == wPos ? _GEN_32 : _GEN_2104;
  assign _GEN_2170 = 6'h17 == wPos ? _GEN_32 : _GEN_2105;
  assign _GEN_2171 = 6'h18 == wPos ? _GEN_32 : _GEN_2106;
  assign _GEN_2172 = 6'h19 == wPos ? _GEN_32 : _GEN_2107;
  assign _GEN_2173 = 6'h1a == wPos ? _GEN_32 : _GEN_2108;
  assign _GEN_2174 = 6'h1b == wPos ? _GEN_32 : _GEN_2109;
  assign _GEN_2175 = 6'h1c == wPos ? _GEN_32 : _GEN_2110;
  assign _GEN_2176 = 6'h1d == wPos ? _GEN_32 : _GEN_2111;
  assign _GEN_2177 = 6'h1e == wPos ? _GEN_32 : _GEN_2112;
  assign _GEN_2178 = 6'h1f == wPos ? _GEN_32 : _GEN_2113;
  assign _GEN_2179 = 6'h20 == wPos ? _GEN_32 : _GEN_2114;
  assign _GEN_2180 = 6'h21 == wPos ? _GEN_32 : _GEN_2115;
  assign _GEN_2181 = 6'h22 == wPos ? _GEN_32 : _GEN_2116;
  assign _GEN_2182 = 6'h23 == wPos ? _GEN_32 : _GEN_2117;
  assign _GEN_2183 = 6'h24 == wPos ? _GEN_32 : _GEN_2118;
  assign _GEN_2184 = 6'h25 == wPos ? _GEN_32 : _GEN_2119;
  assign _GEN_2185 = 6'h26 == wPos ? _GEN_32 : _GEN_2120;
  assign _GEN_2186 = 6'h27 == wPos ? _GEN_32 : _GEN_2121;
  assign _GEN_2187 = 6'h28 == wPos ? _GEN_32 : _GEN_2122;
  assign _GEN_2188 = 6'h29 == wPos ? _GEN_32 : _GEN_2123;
  assign _GEN_2189 = 6'h2a == wPos ? _GEN_32 : _GEN_2124;
  assign _GEN_2190 = 6'h2b == wPos ? _GEN_32 : _GEN_2125;
  assign _GEN_2191 = 6'h2c == wPos ? _GEN_32 : _GEN_2126;
  assign _GEN_2192 = 6'h2d == wPos ? _GEN_32 : _GEN_2127;
  assign _GEN_2193 = 6'h2e == wPos ? _GEN_32 : _GEN_2128;
  assign _GEN_2194 = 6'h2f == wPos ? _GEN_32 : _GEN_2129;
  assign _GEN_2195 = 6'h30 == wPos ? _GEN_32 : _GEN_2130;
  assign _GEN_2196 = 6'h31 == wPos ? _GEN_32 : _GEN_2131;
  assign _GEN_2197 = 6'h32 == wPos ? _GEN_32 : _GEN_2132;
  assign _GEN_2198 = 6'h33 == wPos ? _GEN_32 : _GEN_2133;
  assign _GEN_2199 = 6'h34 == wPos ? _GEN_32 : _GEN_2134;
  assign _GEN_2200 = 6'h35 == wPos ? _GEN_32 : _GEN_2135;
  assign _GEN_2201 = 6'h36 == wPos ? _GEN_32 : _GEN_2136;
  assign _GEN_2202 = 6'h37 == wPos ? _GEN_32 : _GEN_2137;
  assign _GEN_2203 = 6'h38 == wPos ? _GEN_32 : _GEN_2138;
  assign _GEN_2204 = 6'h39 == wPos ? _GEN_32 : _GEN_2139;
  assign _GEN_2205 = 6'h3a == wPos ? _GEN_32 : _GEN_2140;
  assign _GEN_2206 = 6'h3b == wPos ? _GEN_32 : _GEN_2141;
  assign _GEN_2207 = 6'h3c == wPos ? _GEN_32 : _GEN_2142;
  assign _GEN_2208 = 6'h3d == wPos ? _GEN_32 : _GEN_2143;
  assign _GEN_2209 = 6'h3e == wPos ? _GEN_32 : _GEN_2144;
  assign _GEN_2210 = 6'h3f == wPos ? _GEN_32 : _GEN_2145;
  assign _GEN_2211 = _T_149 ? _GEN_2147 : _GEN_2082;
  assign _GEN_2212 = _T_149 ? _GEN_2148 : _GEN_2083;
  assign _GEN_2213 = _T_149 ? _GEN_2149 : _GEN_2084;
  assign _GEN_2214 = _T_149 ? _GEN_2150 : _GEN_2085;
  assign _GEN_2215 = _T_149 ? _GEN_2151 : _GEN_2086;
  assign _GEN_2216 = _T_149 ? _GEN_2152 : _GEN_2087;
  assign _GEN_2217 = _T_149 ? _GEN_2153 : _GEN_2088;
  assign _GEN_2218 = _T_149 ? _GEN_2154 : _GEN_2089;
  assign _GEN_2219 = _T_149 ? _GEN_2155 : _GEN_2090;
  assign _GEN_2220 = _T_149 ? _GEN_2156 : _GEN_2091;
  assign _GEN_2221 = _T_149 ? _GEN_2157 : _GEN_2092;
  assign _GEN_2222 = _T_149 ? _GEN_2158 : _GEN_2093;
  assign _GEN_2223 = _T_149 ? _GEN_2159 : _GEN_2094;
  assign _GEN_2224 = _T_149 ? _GEN_2160 : _GEN_2095;
  assign _GEN_2225 = _T_149 ? _GEN_2161 : _GEN_2096;
  assign _GEN_2226 = _T_149 ? _GEN_2162 : _GEN_2097;
  assign _GEN_2227 = _T_149 ? _GEN_2163 : _GEN_2098;
  assign _GEN_2228 = _T_149 ? _GEN_2164 : _GEN_2099;
  assign _GEN_2229 = _T_149 ? _GEN_2165 : _GEN_2100;
  assign _GEN_2230 = _T_149 ? _GEN_2166 : _GEN_2101;
  assign _GEN_2231 = _T_149 ? _GEN_2167 : _GEN_2102;
  assign _GEN_2232 = _T_149 ? _GEN_2168 : _GEN_2103;
  assign _GEN_2233 = _T_149 ? _GEN_2169 : _GEN_2104;
  assign _GEN_2234 = _T_149 ? _GEN_2170 : _GEN_2105;
  assign _GEN_2235 = _T_149 ? _GEN_2171 : _GEN_2106;
  assign _GEN_2236 = _T_149 ? _GEN_2172 : _GEN_2107;
  assign _GEN_2237 = _T_149 ? _GEN_2173 : _GEN_2108;
  assign _GEN_2238 = _T_149 ? _GEN_2174 : _GEN_2109;
  assign _GEN_2239 = _T_149 ? _GEN_2175 : _GEN_2110;
  assign _GEN_2240 = _T_149 ? _GEN_2176 : _GEN_2111;
  assign _GEN_2241 = _T_149 ? _GEN_2177 : _GEN_2112;
  assign _GEN_2242 = _T_149 ? _GEN_2178 : _GEN_2113;
  assign _GEN_2243 = _T_149 ? _GEN_2179 : _GEN_2114;
  assign _GEN_2244 = _T_149 ? _GEN_2180 : _GEN_2115;
  assign _GEN_2245 = _T_149 ? _GEN_2181 : _GEN_2116;
  assign _GEN_2246 = _T_149 ? _GEN_2182 : _GEN_2117;
  assign _GEN_2247 = _T_149 ? _GEN_2183 : _GEN_2118;
  assign _GEN_2248 = _T_149 ? _GEN_2184 : _GEN_2119;
  assign _GEN_2249 = _T_149 ? _GEN_2185 : _GEN_2120;
  assign _GEN_2250 = _T_149 ? _GEN_2186 : _GEN_2121;
  assign _GEN_2251 = _T_149 ? _GEN_2187 : _GEN_2122;
  assign _GEN_2252 = _T_149 ? _GEN_2188 : _GEN_2123;
  assign _GEN_2253 = _T_149 ? _GEN_2189 : _GEN_2124;
  assign _GEN_2254 = _T_149 ? _GEN_2190 : _GEN_2125;
  assign _GEN_2255 = _T_149 ? _GEN_2191 : _GEN_2126;
  assign _GEN_2256 = _T_149 ? _GEN_2192 : _GEN_2127;
  assign _GEN_2257 = _T_149 ? _GEN_2193 : _GEN_2128;
  assign _GEN_2258 = _T_149 ? _GEN_2194 : _GEN_2129;
  assign _GEN_2259 = _T_149 ? _GEN_2195 : _GEN_2130;
  assign _GEN_2260 = _T_149 ? _GEN_2196 : _GEN_2131;
  assign _GEN_2261 = _T_149 ? _GEN_2197 : _GEN_2132;
  assign _GEN_2262 = _T_149 ? _GEN_2198 : _GEN_2133;
  assign _GEN_2263 = _T_149 ? _GEN_2199 : _GEN_2134;
  assign _GEN_2264 = _T_149 ? _GEN_2200 : _GEN_2135;
  assign _GEN_2265 = _T_149 ? _GEN_2201 : _GEN_2136;
  assign _GEN_2266 = _T_149 ? _GEN_2202 : _GEN_2137;
  assign _GEN_2267 = _T_149 ? _GEN_2203 : _GEN_2138;
  assign _GEN_2268 = _T_149 ? _GEN_2204 : _GEN_2139;
  assign _GEN_2269 = _T_149 ? _GEN_2205 : _GEN_2140;
  assign _GEN_2270 = _T_149 ? _GEN_2206 : _GEN_2141;
  assign _GEN_2271 = _T_149 ? _GEN_2207 : _GEN_2142;
  assign _GEN_2272 = _T_149 ? _GEN_2208 : _GEN_2143;
  assign _GEN_2273 = _T_149 ? _GEN_2209 : _GEN_2144;
  assign _GEN_2274 = _T_149 ? _GEN_2210 : _GEN_2145;
  assign _GEN_2275 = _T_149 ? _T_158 : _GEN_2146;
  assign _T_323 = _T_149 == 1'h0;
  assign _GEN_2276 = _T_323 ? io_in : _GEN_2211;
  assign _GEN_2277 = _T_323 ? 6'h1 : _GEN_2275;
  assign _GEN_2278 = _T_323 ? 3'h0 : rPos;
  assign _GEN_2279 = io_push ? _GEN_2276 : _GEN_2082;
  assign _GEN_2280 = io_push ? _GEN_2212 : _GEN_2083;
  assign _GEN_2281 = io_push ? _GEN_2213 : _GEN_2084;
  assign _GEN_2282 = io_push ? _GEN_2214 : _GEN_2085;
  assign _GEN_2283 = io_push ? _GEN_2215 : _GEN_2086;
  assign _GEN_2284 = io_push ? _GEN_2216 : _GEN_2087;
  assign _GEN_2285 = io_push ? _GEN_2217 : _GEN_2088;
  assign _GEN_2286 = io_push ? _GEN_2218 : _GEN_2089;
  assign _GEN_2287 = io_push ? _GEN_2219 : _GEN_2090;
  assign _GEN_2288 = io_push ? _GEN_2220 : _GEN_2091;
  assign _GEN_2289 = io_push ? _GEN_2221 : _GEN_2092;
  assign _GEN_2290 = io_push ? _GEN_2222 : _GEN_2093;
  assign _GEN_2291 = io_push ? _GEN_2223 : _GEN_2094;
  assign _GEN_2292 = io_push ? _GEN_2224 : _GEN_2095;
  assign _GEN_2293 = io_push ? _GEN_2225 : _GEN_2096;
  assign _GEN_2294 = io_push ? _GEN_2226 : _GEN_2097;
  assign _GEN_2295 = io_push ? _GEN_2227 : _GEN_2098;
  assign _GEN_2296 = io_push ? _GEN_2228 : _GEN_2099;
  assign _GEN_2297 = io_push ? _GEN_2229 : _GEN_2100;
  assign _GEN_2298 = io_push ? _GEN_2230 : _GEN_2101;
  assign _GEN_2299 = io_push ? _GEN_2231 : _GEN_2102;
  assign _GEN_2300 = io_push ? _GEN_2232 : _GEN_2103;
  assign _GEN_2301 = io_push ? _GEN_2233 : _GEN_2104;
  assign _GEN_2302 = io_push ? _GEN_2234 : _GEN_2105;
  assign _GEN_2303 = io_push ? _GEN_2235 : _GEN_2106;
  assign _GEN_2304 = io_push ? _GEN_2236 : _GEN_2107;
  assign _GEN_2305 = io_push ? _GEN_2237 : _GEN_2108;
  assign _GEN_2306 = io_push ? _GEN_2238 : _GEN_2109;
  assign _GEN_2307 = io_push ? _GEN_2239 : _GEN_2110;
  assign _GEN_2308 = io_push ? _GEN_2240 : _GEN_2111;
  assign _GEN_2309 = io_push ? _GEN_2241 : _GEN_2112;
  assign _GEN_2310 = io_push ? _GEN_2242 : _GEN_2113;
  assign _GEN_2311 = io_push ? _GEN_2243 : _GEN_2114;
  assign _GEN_2312 = io_push ? _GEN_2244 : _GEN_2115;
  assign _GEN_2313 = io_push ? _GEN_2245 : _GEN_2116;
  assign _GEN_2314 = io_push ? _GEN_2246 : _GEN_2117;
  assign _GEN_2315 = io_push ? _GEN_2247 : _GEN_2118;
  assign _GEN_2316 = io_push ? _GEN_2248 : _GEN_2119;
  assign _GEN_2317 = io_push ? _GEN_2249 : _GEN_2120;
  assign _GEN_2318 = io_push ? _GEN_2250 : _GEN_2121;
  assign _GEN_2319 = io_push ? _GEN_2251 : _GEN_2122;
  assign _GEN_2320 = io_push ? _GEN_2252 : _GEN_2123;
  assign _GEN_2321 = io_push ? _GEN_2253 : _GEN_2124;
  assign _GEN_2322 = io_push ? _GEN_2254 : _GEN_2125;
  assign _GEN_2323 = io_push ? _GEN_2255 : _GEN_2126;
  assign _GEN_2324 = io_push ? _GEN_2256 : _GEN_2127;
  assign _GEN_2325 = io_push ? _GEN_2257 : _GEN_2128;
  assign _GEN_2326 = io_push ? _GEN_2258 : _GEN_2129;
  assign _GEN_2327 = io_push ? _GEN_2259 : _GEN_2130;
  assign _GEN_2328 = io_push ? _GEN_2260 : _GEN_2131;
  assign _GEN_2329 = io_push ? _GEN_2261 : _GEN_2132;
  assign _GEN_2330 = io_push ? _GEN_2262 : _GEN_2133;
  assign _GEN_2331 = io_push ? _GEN_2263 : _GEN_2134;
  assign _GEN_2332 = io_push ? _GEN_2264 : _GEN_2135;
  assign _GEN_2333 = io_push ? _GEN_2265 : _GEN_2136;
  assign _GEN_2334 = io_push ? _GEN_2266 : _GEN_2137;
  assign _GEN_2335 = io_push ? _GEN_2267 : _GEN_2138;
  assign _GEN_2336 = io_push ? _GEN_2268 : _GEN_2139;
  assign _GEN_2337 = io_push ? _GEN_2269 : _GEN_2140;
  assign _GEN_2338 = io_push ? _GEN_2270 : _GEN_2141;
  assign _GEN_2339 = io_push ? _GEN_2271 : _GEN_2142;
  assign _GEN_2340 = io_push ? _GEN_2272 : _GEN_2143;
  assign _GEN_2341 = io_push ? _GEN_2273 : _GEN_2144;
  assign _GEN_2342 = io_push ? _GEN_2274 : _GEN_2145;
  assign _GEN_2343 = io_push ? _GEN_2277 : _GEN_2146;
  assign _GEN_2344 = io_push ? _GEN_2278 : rPos;
  assign _T_329 = rPos + 3'h1;
  assign _T_330 = _T_329[2:0];
  assign _GEN_2345 = _T_149 ? _T_330 : _GEN_2344;
  assign _GEN_2346 = _T_323 ? 3'h1 : _GEN_2345;
  assign _GEN_2347 = _T_323 ? 6'h0 : _GEN_2343;
  assign _GEN_2348 = io_pop ? _GEN_2346 : _GEN_2344;
  assign _GEN_2349 = io_pop ? _GEN_2347 : _GEN_2343;
  assign _GEN_2350 = _T_315 ? _GEN_2279 : _GEN_2082;
  assign _GEN_2351 = _T_315 ? _GEN_2280 : _GEN_2083;
  assign _GEN_2352 = _T_315 ? _GEN_2281 : _GEN_2084;
  assign _GEN_2353 = _T_315 ? _GEN_2282 : _GEN_2085;
  assign _GEN_2354 = _T_315 ? _GEN_2283 : _GEN_2086;
  assign _GEN_2355 = _T_315 ? _GEN_2284 : _GEN_2087;
  assign _GEN_2356 = _T_315 ? _GEN_2285 : _GEN_2088;
  assign _GEN_2357 = _T_315 ? _GEN_2286 : _GEN_2089;
  assign _GEN_2358 = _T_315 ? _GEN_2287 : _GEN_2090;
  assign _GEN_2359 = _T_315 ? _GEN_2288 : _GEN_2091;
  assign _GEN_2360 = _T_315 ? _GEN_2289 : _GEN_2092;
  assign _GEN_2361 = _T_315 ? _GEN_2290 : _GEN_2093;
  assign _GEN_2362 = _T_315 ? _GEN_2291 : _GEN_2094;
  assign _GEN_2363 = _T_315 ? _GEN_2292 : _GEN_2095;
  assign _GEN_2364 = _T_315 ? _GEN_2293 : _GEN_2096;
  assign _GEN_2365 = _T_315 ? _GEN_2294 : _GEN_2097;
  assign _GEN_2366 = _T_315 ? _GEN_2295 : _GEN_2098;
  assign _GEN_2367 = _T_315 ? _GEN_2296 : _GEN_2099;
  assign _GEN_2368 = _T_315 ? _GEN_2297 : _GEN_2100;
  assign _GEN_2369 = _T_315 ? _GEN_2298 : _GEN_2101;
  assign _GEN_2370 = _T_315 ? _GEN_2299 : _GEN_2102;
  assign _GEN_2371 = _T_315 ? _GEN_2300 : _GEN_2103;
  assign _GEN_2372 = _T_315 ? _GEN_2301 : _GEN_2104;
  assign _GEN_2373 = _T_315 ? _GEN_2302 : _GEN_2105;
  assign _GEN_2374 = _T_315 ? _GEN_2303 : _GEN_2106;
  assign _GEN_2375 = _T_315 ? _GEN_2304 : _GEN_2107;
  assign _GEN_2376 = _T_315 ? _GEN_2305 : _GEN_2108;
  assign _GEN_2377 = _T_315 ? _GEN_2306 : _GEN_2109;
  assign _GEN_2378 = _T_315 ? _GEN_2307 : _GEN_2110;
  assign _GEN_2379 = _T_315 ? _GEN_2308 : _GEN_2111;
  assign _GEN_2380 = _T_315 ? _GEN_2309 : _GEN_2112;
  assign _GEN_2381 = _T_315 ? _GEN_2310 : _GEN_2113;
  assign _GEN_2382 = _T_315 ? _GEN_2311 : _GEN_2114;
  assign _GEN_2383 = _T_315 ? _GEN_2312 : _GEN_2115;
  assign _GEN_2384 = _T_315 ? _GEN_2313 : _GEN_2116;
  assign _GEN_2385 = _T_315 ? _GEN_2314 : _GEN_2117;
  assign _GEN_2386 = _T_315 ? _GEN_2315 : _GEN_2118;
  assign _GEN_2387 = _T_315 ? _GEN_2316 : _GEN_2119;
  assign _GEN_2388 = _T_315 ? _GEN_2317 : _GEN_2120;
  assign _GEN_2389 = _T_315 ? _GEN_2318 : _GEN_2121;
  assign _GEN_2390 = _T_315 ? _GEN_2319 : _GEN_2122;
  assign _GEN_2391 = _T_315 ? _GEN_2320 : _GEN_2123;
  assign _GEN_2392 = _T_315 ? _GEN_2321 : _GEN_2124;
  assign _GEN_2393 = _T_315 ? _GEN_2322 : _GEN_2125;
  assign _GEN_2394 = _T_315 ? _GEN_2323 : _GEN_2126;
  assign _GEN_2395 = _T_315 ? _GEN_2324 : _GEN_2127;
  assign _GEN_2396 = _T_315 ? _GEN_2325 : _GEN_2128;
  assign _GEN_2397 = _T_315 ? _GEN_2326 : _GEN_2129;
  assign _GEN_2398 = _T_315 ? _GEN_2327 : _GEN_2130;
  assign _GEN_2399 = _T_315 ? _GEN_2328 : _GEN_2131;
  assign _GEN_2400 = _T_315 ? _GEN_2329 : _GEN_2132;
  assign _GEN_2401 = _T_315 ? _GEN_2330 : _GEN_2133;
  assign _GEN_2402 = _T_315 ? _GEN_2331 : _GEN_2134;
  assign _GEN_2403 = _T_315 ? _GEN_2332 : _GEN_2135;
  assign _GEN_2404 = _T_315 ? _GEN_2333 : _GEN_2136;
  assign _GEN_2405 = _T_315 ? _GEN_2334 : _GEN_2137;
  assign _GEN_2406 = _T_315 ? _GEN_2335 : _GEN_2138;
  assign _GEN_2407 = _T_315 ? _GEN_2336 : _GEN_2139;
  assign _GEN_2408 = _T_315 ? _GEN_2337 : _GEN_2140;
  assign _GEN_2409 = _T_315 ? _GEN_2338 : _GEN_2141;
  assign _GEN_2410 = _T_315 ? _GEN_2339 : _GEN_2142;
  assign _GEN_2411 = _T_315 ? _GEN_2340 : _GEN_2143;
  assign _GEN_2412 = _T_315 ? _GEN_2341 : _GEN_2144;
  assign _GEN_2413 = _T_315 ? _GEN_2342 : _GEN_2145;
  assign _GEN_2414 = _T_315 ? _GEN_2349 : _GEN_2146;
  assign _GEN_2415 = _T_315 ? _GEN_2348 : rPos;
  assign _T_336 = io_pop == 1'h0;
  assign _T_337 = io_reset & _T_336;
  assign _T_339 = io_push == 1'h0;
  assign _T_340 = _T_337 & _T_339;
  assign _GEN_2416 = _T_340 ? 6'h0 : _GEN_2414;
  assign _GEN_2417 = _T_340 ? 3'h0 : _GEN_2415;
  assign _GEN_33 = _GEN_2424;
  assign _GEN_2418 = 3'h1 == rPos ? catMem_1 : catMem_0;
  assign _GEN_2419 = 3'h2 == rPos ? catMem_2 : _GEN_2418;
  assign _GEN_2420 = 3'h3 == rPos ? catMem_3 : _GEN_2419;
  assign _GEN_2421 = 3'h4 == rPos ? catMem_4 : _GEN_2420;
  assign _GEN_2422 = 3'h5 == rPos ? catMem_5 : _GEN_2421;
  assign _GEN_2423 = 3'h6 == rPos ? catMem_6 : _GEN_2422;
  assign _GEN_2424 = 3'h7 == rPos ? catMem_7 : _GEN_2423;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2425 = {1{$random}};
  wPos = _GEN_2425[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2426 = {1{$random}};
  rPos = _GEN_2426[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2427 = {1{$random}};
  mem_0 = _GEN_2427[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2428 = {1{$random}};
  mem_1 = _GEN_2428[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2429 = {1{$random}};
  mem_2 = _GEN_2429[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2430 = {1{$random}};
  mem_3 = _GEN_2430[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2431 = {1{$random}};
  mem_4 = _GEN_2431[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2432 = {1{$random}};
  mem_5 = _GEN_2432[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2433 = {1{$random}};
  mem_6 = _GEN_2433[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2434 = {1{$random}};
  mem_7 = _GEN_2434[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2435 = {1{$random}};
  mem_8 = _GEN_2435[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2436 = {1{$random}};
  mem_9 = _GEN_2436[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2437 = {1{$random}};
  mem_10 = _GEN_2437[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2438 = {1{$random}};
  mem_11 = _GEN_2438[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2439 = {1{$random}};
  mem_12 = _GEN_2439[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2440 = {1{$random}};
  mem_13 = _GEN_2440[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2441 = {1{$random}};
  mem_14 = _GEN_2441[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2442 = {1{$random}};
  mem_15 = _GEN_2442[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2443 = {1{$random}};
  mem_16 = _GEN_2443[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2444 = {1{$random}};
  mem_17 = _GEN_2444[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2445 = {1{$random}};
  mem_18 = _GEN_2445[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2446 = {1{$random}};
  mem_19 = _GEN_2446[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2447 = {1{$random}};
  mem_20 = _GEN_2447[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2448 = {1{$random}};
  mem_21 = _GEN_2448[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2449 = {1{$random}};
  mem_22 = _GEN_2449[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2450 = {1{$random}};
  mem_23 = _GEN_2450[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2451 = {1{$random}};
  mem_24 = _GEN_2451[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2452 = {1{$random}};
  mem_25 = _GEN_2452[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2453 = {1{$random}};
  mem_26 = _GEN_2453[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2454 = {1{$random}};
  mem_27 = _GEN_2454[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2455 = {1{$random}};
  mem_28 = _GEN_2455[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2456 = {1{$random}};
  mem_29 = _GEN_2456[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2457 = {1{$random}};
  mem_30 = _GEN_2457[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2458 = {1{$random}};
  mem_31 = _GEN_2458[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2459 = {1{$random}};
  mem_32 = _GEN_2459[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2460 = {1{$random}};
  mem_33 = _GEN_2460[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2461 = {1{$random}};
  mem_34 = _GEN_2461[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2462 = {1{$random}};
  mem_35 = _GEN_2462[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2463 = {1{$random}};
  mem_36 = _GEN_2463[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2464 = {1{$random}};
  mem_37 = _GEN_2464[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2465 = {1{$random}};
  mem_38 = _GEN_2465[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2466 = {1{$random}};
  mem_39 = _GEN_2466[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2467 = {1{$random}};
  mem_40 = _GEN_2467[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2468 = {1{$random}};
  mem_41 = _GEN_2468[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2469 = {1{$random}};
  mem_42 = _GEN_2469[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2470 = {1{$random}};
  mem_43 = _GEN_2470[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2471 = {1{$random}};
  mem_44 = _GEN_2471[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2472 = {1{$random}};
  mem_45 = _GEN_2472[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2473 = {1{$random}};
  mem_46 = _GEN_2473[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2474 = {1{$random}};
  mem_47 = _GEN_2474[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2475 = {1{$random}};
  mem_48 = _GEN_2475[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2476 = {1{$random}};
  mem_49 = _GEN_2476[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2477 = {1{$random}};
  mem_50 = _GEN_2477[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2478 = {1{$random}};
  mem_51 = _GEN_2478[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2479 = {1{$random}};
  mem_52 = _GEN_2479[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2480 = {1{$random}};
  mem_53 = _GEN_2480[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2481 = {1{$random}};
  mem_54 = _GEN_2481[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2482 = {1{$random}};
  mem_55 = _GEN_2482[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2483 = {1{$random}};
  mem_56 = _GEN_2483[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2484 = {1{$random}};
  mem_57 = _GEN_2484[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2485 = {1{$random}};
  mem_58 = _GEN_2485[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2486 = {1{$random}};
  mem_59 = _GEN_2486[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2487 = {1{$random}};
  mem_60 = _GEN_2487[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2488 = {1{$random}};
  mem_61 = _GEN_2488[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2489 = {1{$random}};
  mem_62 = _GEN_2489[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2490 = {1{$random}};
  mem_63 = _GEN_2490[3:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (_T_340) begin
      wPos <= 6'h0;
    end else begin
      if (_T_315) begin
        if (io_pop) begin
          if (_T_323) begin
            wPos <= 6'h0;
          end else begin
            if (io_push) begin
              if (_T_323) begin
                wPos <= 6'h1;
              end else begin
                if (_T_149) begin
                  wPos <= _T_158;
                end else begin
                  if (_T_150) begin
                    wPos <= _T_313;
                  end
                end
              end
            end else begin
              if (_T_150) begin
                wPos <= _T_313;
              end
            end
          end
        end else begin
          if (io_push) begin
            if (_T_323) begin
              wPos <= 6'h1;
            end else begin
              if (_T_149) begin
                wPos <= _T_158;
              end else begin
                if (_T_150) begin
                  wPos <= _T_313;
                end
              end
            end
          end else begin
            if (_T_150) begin
              wPos <= _T_313;
            end
          end
        end
      end else begin
        wPos <= _GEN_2146;
      end
    end
    if (_T_340) begin
      rPos <= 3'h0;
    end else begin
      if (_T_315) begin
        if (io_pop) begin
          if (_T_323) begin
            rPos <= 3'h1;
          end else begin
            if (_T_149) begin
              rPos <= _T_330;
            end else begin
              if (io_push) begin
                if (_T_323) begin
                  rPos <= 3'h0;
                end
              end
            end
          end
        end else begin
          if (io_push) begin
            if (_T_323) begin
              rPos <= 3'h0;
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_323) begin
          mem_0 <= io_in;
        end else begin
          if (_T_149) begin
            if (6'h0 == wPos) begin
              mem_0 <= _GEN_32;
            end else begin
              if (_T_150) begin
                if (6'h0 == _T_308) begin
                  mem_0 <= _GEN_31;
                end else begin
                  if (6'h0 == _T_303) begin
                    mem_0 <= _GEN_30;
                  end else begin
                    if (6'h0 == _T_298) begin
                      mem_0 <= _GEN_29;
                    end else begin
                      if (6'h0 == _T_293) begin
                        mem_0 <= _GEN_28;
                      end else begin
                        if (6'h0 == _T_288) begin
                          mem_0 <= _GEN_27;
                        end else begin
                          if (6'h0 == _T_283) begin
                            mem_0 <= _GEN_26;
                          end else begin
                            if (6'h0 == _T_278) begin
                              mem_0 <= _GEN_25;
                            end else begin
                              if (6'h0 == _T_273) begin
                                mem_0 <= _GEN_24;
                              end else begin
                                if (6'h0 == _T_268) begin
                                  mem_0 <= _GEN_23;
                                end else begin
                                  if (6'h0 == _T_263) begin
                                    mem_0 <= _GEN_22;
                                  end else begin
                                    if (6'h0 == _T_258) begin
                                      mem_0 <= _GEN_21;
                                    end else begin
                                      if (6'h0 == _T_253) begin
                                        mem_0 <= _GEN_20;
                                      end else begin
                                        if (6'h0 == _T_248) begin
                                          mem_0 <= _GEN_19;
                                        end else begin
                                          if (6'h0 == _T_243) begin
                                            mem_0 <= _GEN_18;
                                          end else begin
                                            if (6'h0 == _T_238) begin
                                              mem_0 <= _GEN_17;
                                            end else begin
                                              if (6'h0 == _T_233) begin
                                                mem_0 <= _GEN_16;
                                              end else begin
                                                if (6'h0 == _T_228) begin
                                                  mem_0 <= _GEN_15;
                                                end else begin
                                                  if (6'h0 == _T_223) begin
                                                    mem_0 <= _GEN_14;
                                                  end else begin
                                                    if (6'h0 == _T_218) begin
                                                      mem_0 <= _GEN_13;
                                                    end else begin
                                                      if (6'h0 == _T_213) begin
                                                        mem_0 <= _GEN_12;
                                                      end else begin
                                                        if (6'h0 == _T_208) begin
                                                          mem_0 <= _GEN_11;
                                                        end else begin
                                                          if (6'h0 == _T_203) begin
                                                            mem_0 <= _GEN_10;
                                                          end else begin
                                                            if (6'h0 == _T_198) begin
                                                              mem_0 <= _GEN_9;
                                                            end else begin
                                                              if (6'h0 == _T_193) begin
                                                                mem_0 <= _GEN_8;
                                                              end else begin
                                                                if (6'h0 == _T_188) begin
                                                                  mem_0 <= _GEN_7;
                                                                end else begin
                                                                  if (6'h0 == _T_183) begin
                                                                    mem_0 <= _GEN_6;
                                                                  end else begin
                                                                    if (6'h0 == _T_178) begin
                                                                      mem_0 <= _GEN_5;
                                                                    end else begin
                                                                      if (6'h0 == _T_173) begin
                                                                        mem_0 <= _GEN_4;
                                                                      end else begin
                                                                        if (6'h0 == _T_168) begin
                                                                          mem_0 <= _GEN_3;
                                                                        end else begin
                                                                          if (6'h0 == _T_163) begin
                                                                            mem_0 <= _GEN_2;
                                                                          end else begin
                                                                            if (6'h0 == _T_158) begin
                                                                              mem_0 <= _GEN_1;
                                                                            end else begin
                                                                              if (6'h0 == _T_153) begin
                                                                                mem_0 <= _GEN_0;
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_150) begin
              if (6'h0 == _T_308) begin
                mem_0 <= _GEN_31;
              end else begin
                if (6'h0 == _T_303) begin
                  mem_0 <= _GEN_30;
                end else begin
                  if (6'h0 == _T_298) begin
                    mem_0 <= _GEN_29;
                  end else begin
                    if (6'h0 == _T_293) begin
                      mem_0 <= _GEN_28;
                    end else begin
                      if (6'h0 == _T_288) begin
                        mem_0 <= _GEN_27;
                      end else begin
                        if (6'h0 == _T_283) begin
                          mem_0 <= _GEN_26;
                        end else begin
                          if (6'h0 == _T_278) begin
                            mem_0 <= _GEN_25;
                          end else begin
                            if (6'h0 == _T_273) begin
                              mem_0 <= _GEN_24;
                            end else begin
                              if (6'h0 == _T_268) begin
                                mem_0 <= _GEN_23;
                              end else begin
                                if (6'h0 == _T_263) begin
                                  mem_0 <= _GEN_22;
                                end else begin
                                  if (6'h0 == _T_258) begin
                                    mem_0 <= _GEN_21;
                                  end else begin
                                    if (6'h0 == _T_253) begin
                                      mem_0 <= _GEN_20;
                                    end else begin
                                      if (6'h0 == _T_248) begin
                                        mem_0 <= _GEN_19;
                                      end else begin
                                        if (6'h0 == _T_243) begin
                                          mem_0 <= _GEN_18;
                                        end else begin
                                          if (6'h0 == _T_238) begin
                                            mem_0 <= _GEN_17;
                                          end else begin
                                            if (6'h0 == _T_233) begin
                                              mem_0 <= _GEN_16;
                                            end else begin
                                              if (6'h0 == _T_228) begin
                                                mem_0 <= _GEN_15;
                                              end else begin
                                                if (6'h0 == _T_223) begin
                                                  mem_0 <= _GEN_14;
                                                end else begin
                                                  if (6'h0 == _T_218) begin
                                                    mem_0 <= _GEN_13;
                                                  end else begin
                                                    if (6'h0 == _T_213) begin
                                                      mem_0 <= _GEN_12;
                                                    end else begin
                                                      if (6'h0 == _T_208) begin
                                                        mem_0 <= _GEN_11;
                                                      end else begin
                                                        if (6'h0 == _T_203) begin
                                                          mem_0 <= _GEN_10;
                                                        end else begin
                                                          if (6'h0 == _T_198) begin
                                                            mem_0 <= _GEN_9;
                                                          end else begin
                                                            if (6'h0 == _T_193) begin
                                                              mem_0 <= _GEN_8;
                                                            end else begin
                                                              if (6'h0 == _T_188) begin
                                                                mem_0 <= _GEN_7;
                                                              end else begin
                                                                if (6'h0 == _T_183) begin
                                                                  mem_0 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h0 == _T_178) begin
                                                                    mem_0 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h0 == _T_173) begin
                                                                      mem_0 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h0 == _T_168) begin
                                                                        mem_0 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h0 == _T_163) begin
                                                                          mem_0 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h0 == _T_158) begin
                                                                            mem_0 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h0 == _T_153) begin
                                                                              mem_0 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h0 == _T_308) begin
            mem_0 <= _GEN_31;
          end else begin
            if (6'h0 == _T_303) begin
              mem_0 <= _GEN_30;
            end else begin
              if (6'h0 == _T_298) begin
                mem_0 <= _GEN_29;
              end else begin
                if (6'h0 == _T_293) begin
                  mem_0 <= _GEN_28;
                end else begin
                  if (6'h0 == _T_288) begin
                    mem_0 <= _GEN_27;
                  end else begin
                    if (6'h0 == _T_283) begin
                      mem_0 <= _GEN_26;
                    end else begin
                      if (6'h0 == _T_278) begin
                        mem_0 <= _GEN_25;
                      end else begin
                        if (6'h0 == _T_273) begin
                          mem_0 <= _GEN_24;
                        end else begin
                          if (6'h0 == _T_268) begin
                            mem_0 <= _GEN_23;
                          end else begin
                            if (6'h0 == _T_263) begin
                              mem_0 <= _GEN_22;
                            end else begin
                              if (6'h0 == _T_258) begin
                                mem_0 <= _GEN_21;
                              end else begin
                                if (6'h0 == _T_253) begin
                                  mem_0 <= _GEN_20;
                                end else begin
                                  if (6'h0 == _T_248) begin
                                    mem_0 <= _GEN_19;
                                  end else begin
                                    if (6'h0 == _T_243) begin
                                      mem_0 <= _GEN_18;
                                    end else begin
                                      if (6'h0 == _T_238) begin
                                        mem_0 <= _GEN_17;
                                      end else begin
                                        if (6'h0 == _T_233) begin
                                          mem_0 <= _GEN_16;
                                        end else begin
                                          if (6'h0 == _T_228) begin
                                            mem_0 <= _GEN_15;
                                          end else begin
                                            if (6'h0 == _T_223) begin
                                              mem_0 <= _GEN_14;
                                            end else begin
                                              if (6'h0 == _T_218) begin
                                                mem_0 <= _GEN_13;
                                              end else begin
                                                if (6'h0 == _T_213) begin
                                                  mem_0 <= _GEN_12;
                                                end else begin
                                                  if (6'h0 == _T_208) begin
                                                    mem_0 <= _GEN_11;
                                                  end else begin
                                                    if (6'h0 == _T_203) begin
                                                      mem_0 <= _GEN_10;
                                                    end else begin
                                                      if (6'h0 == _T_198) begin
                                                        mem_0 <= _GEN_9;
                                                      end else begin
                                                        if (6'h0 == _T_193) begin
                                                          mem_0 <= _GEN_8;
                                                        end else begin
                                                          if (6'h0 == _T_188) begin
                                                            mem_0 <= _GEN_7;
                                                          end else begin
                                                            if (6'h0 == _T_183) begin
                                                              mem_0 <= _GEN_6;
                                                            end else begin
                                                              if (6'h0 == _T_178) begin
                                                                mem_0 <= _GEN_5;
                                                              end else begin
                                                                if (6'h0 == _T_173) begin
                                                                  mem_0 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h0 == _T_168) begin
                                                                    mem_0 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h0 == _T_163) begin
                                                                      mem_0 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h0 == _T_158) begin
                                                                        mem_0 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h0 == _T_153) begin
                                                                          mem_0 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h0 == _T_308) begin
          mem_0 <= _GEN_31;
        end else begin
          if (6'h0 == _T_303) begin
            mem_0 <= _GEN_30;
          end else begin
            if (6'h0 == _T_298) begin
              mem_0 <= _GEN_29;
            end else begin
              if (6'h0 == _T_293) begin
                mem_0 <= _GEN_28;
              end else begin
                if (6'h0 == _T_288) begin
                  mem_0 <= _GEN_27;
                end else begin
                  if (6'h0 == _T_283) begin
                    mem_0 <= _GEN_26;
                  end else begin
                    if (6'h0 == _T_278) begin
                      mem_0 <= _GEN_25;
                    end else begin
                      if (6'h0 == _T_273) begin
                        mem_0 <= _GEN_24;
                      end else begin
                        if (6'h0 == _T_268) begin
                          mem_0 <= _GEN_23;
                        end else begin
                          if (6'h0 == _T_263) begin
                            mem_0 <= _GEN_22;
                          end else begin
                            if (6'h0 == _T_258) begin
                              mem_0 <= _GEN_21;
                            end else begin
                              if (6'h0 == _T_253) begin
                                mem_0 <= _GEN_20;
                              end else begin
                                if (6'h0 == _T_248) begin
                                  mem_0 <= _GEN_19;
                                end else begin
                                  if (6'h0 == _T_243) begin
                                    mem_0 <= _GEN_18;
                                  end else begin
                                    if (6'h0 == _T_238) begin
                                      mem_0 <= _GEN_17;
                                    end else begin
                                      if (6'h0 == _T_233) begin
                                        mem_0 <= _GEN_16;
                                      end else begin
                                        if (6'h0 == _T_228) begin
                                          mem_0 <= _GEN_15;
                                        end else begin
                                          if (6'h0 == _T_223) begin
                                            mem_0 <= _GEN_14;
                                          end else begin
                                            if (6'h0 == _T_218) begin
                                              mem_0 <= _GEN_13;
                                            end else begin
                                              if (6'h0 == _T_213) begin
                                                mem_0 <= _GEN_12;
                                              end else begin
                                                if (6'h0 == _T_208) begin
                                                  mem_0 <= _GEN_11;
                                                end else begin
                                                  if (6'h0 == _T_203) begin
                                                    mem_0 <= _GEN_10;
                                                  end else begin
                                                    if (6'h0 == _T_198) begin
                                                      mem_0 <= _GEN_9;
                                                    end else begin
                                                      if (6'h0 == _T_193) begin
                                                        mem_0 <= _GEN_8;
                                                      end else begin
                                                        if (6'h0 == _T_188) begin
                                                          mem_0 <= _GEN_7;
                                                        end else begin
                                                          if (6'h0 == _T_183) begin
                                                            mem_0 <= _GEN_6;
                                                          end else begin
                                                            if (6'h0 == _T_178) begin
                                                              mem_0 <= _GEN_5;
                                                            end else begin
                                                              if (6'h0 == _T_173) begin
                                                                mem_0 <= _GEN_4;
                                                              end else begin
                                                                if (6'h0 == _T_168) begin
                                                                  mem_0 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h0 == _T_163) begin
                                                                    mem_0 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h0 == _T_158) begin
                                                                      mem_0 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h0 == _T_153) begin
                                                                        mem_0 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h1 == wPos) begin
            mem_1 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h1 == _T_308) begin
                mem_1 <= _GEN_31;
              end else begin
                if (6'h1 == _T_303) begin
                  mem_1 <= _GEN_30;
                end else begin
                  if (6'h1 == _T_298) begin
                    mem_1 <= _GEN_29;
                  end else begin
                    if (6'h1 == _T_293) begin
                      mem_1 <= _GEN_28;
                    end else begin
                      if (6'h1 == _T_288) begin
                        mem_1 <= _GEN_27;
                      end else begin
                        if (6'h1 == _T_283) begin
                          mem_1 <= _GEN_26;
                        end else begin
                          if (6'h1 == _T_278) begin
                            mem_1 <= _GEN_25;
                          end else begin
                            if (6'h1 == _T_273) begin
                              mem_1 <= _GEN_24;
                            end else begin
                              if (6'h1 == _T_268) begin
                                mem_1 <= _GEN_23;
                              end else begin
                                if (6'h1 == _T_263) begin
                                  mem_1 <= _GEN_22;
                                end else begin
                                  if (6'h1 == _T_258) begin
                                    mem_1 <= _GEN_21;
                                  end else begin
                                    if (6'h1 == _T_253) begin
                                      mem_1 <= _GEN_20;
                                    end else begin
                                      if (6'h1 == _T_248) begin
                                        mem_1 <= _GEN_19;
                                      end else begin
                                        if (6'h1 == _T_243) begin
                                          mem_1 <= _GEN_18;
                                        end else begin
                                          if (6'h1 == _T_238) begin
                                            mem_1 <= _GEN_17;
                                          end else begin
                                            if (6'h1 == _T_233) begin
                                              mem_1 <= _GEN_16;
                                            end else begin
                                              if (6'h1 == _T_228) begin
                                                mem_1 <= _GEN_15;
                                              end else begin
                                                if (6'h1 == _T_223) begin
                                                  mem_1 <= _GEN_14;
                                                end else begin
                                                  if (6'h1 == _T_218) begin
                                                    mem_1 <= _GEN_13;
                                                  end else begin
                                                    if (6'h1 == _T_213) begin
                                                      mem_1 <= _GEN_12;
                                                    end else begin
                                                      if (6'h1 == _T_208) begin
                                                        mem_1 <= _GEN_11;
                                                      end else begin
                                                        if (6'h1 == _T_203) begin
                                                          mem_1 <= _GEN_10;
                                                        end else begin
                                                          if (6'h1 == _T_198) begin
                                                            mem_1 <= _GEN_9;
                                                          end else begin
                                                            if (6'h1 == _T_193) begin
                                                              mem_1 <= _GEN_8;
                                                            end else begin
                                                              if (6'h1 == _T_188) begin
                                                                mem_1 <= _GEN_7;
                                                              end else begin
                                                                if (6'h1 == _T_183) begin
                                                                  mem_1 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h1 == _T_178) begin
                                                                    mem_1 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h1 == _T_173) begin
                                                                      mem_1 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h1 == _T_168) begin
                                                                        mem_1 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h1 == _T_163) begin
                                                                          mem_1 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h1 == _T_158) begin
                                                                            mem_1 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h1 == _T_153) begin
                                                                              mem_1 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h1 == _T_308) begin
              mem_1 <= _GEN_31;
            end else begin
              if (6'h1 == _T_303) begin
                mem_1 <= _GEN_30;
              end else begin
                if (6'h1 == _T_298) begin
                  mem_1 <= _GEN_29;
                end else begin
                  if (6'h1 == _T_293) begin
                    mem_1 <= _GEN_28;
                  end else begin
                    if (6'h1 == _T_288) begin
                      mem_1 <= _GEN_27;
                    end else begin
                      if (6'h1 == _T_283) begin
                        mem_1 <= _GEN_26;
                      end else begin
                        if (6'h1 == _T_278) begin
                          mem_1 <= _GEN_25;
                        end else begin
                          if (6'h1 == _T_273) begin
                            mem_1 <= _GEN_24;
                          end else begin
                            if (6'h1 == _T_268) begin
                              mem_1 <= _GEN_23;
                            end else begin
                              if (6'h1 == _T_263) begin
                                mem_1 <= _GEN_22;
                              end else begin
                                if (6'h1 == _T_258) begin
                                  mem_1 <= _GEN_21;
                                end else begin
                                  if (6'h1 == _T_253) begin
                                    mem_1 <= _GEN_20;
                                  end else begin
                                    if (6'h1 == _T_248) begin
                                      mem_1 <= _GEN_19;
                                    end else begin
                                      if (6'h1 == _T_243) begin
                                        mem_1 <= _GEN_18;
                                      end else begin
                                        if (6'h1 == _T_238) begin
                                          mem_1 <= _GEN_17;
                                        end else begin
                                          if (6'h1 == _T_233) begin
                                            mem_1 <= _GEN_16;
                                          end else begin
                                            if (6'h1 == _T_228) begin
                                              mem_1 <= _GEN_15;
                                            end else begin
                                              if (6'h1 == _T_223) begin
                                                mem_1 <= _GEN_14;
                                              end else begin
                                                if (6'h1 == _T_218) begin
                                                  mem_1 <= _GEN_13;
                                                end else begin
                                                  if (6'h1 == _T_213) begin
                                                    mem_1 <= _GEN_12;
                                                  end else begin
                                                    if (6'h1 == _T_208) begin
                                                      mem_1 <= _GEN_11;
                                                    end else begin
                                                      if (6'h1 == _T_203) begin
                                                        mem_1 <= _GEN_10;
                                                      end else begin
                                                        if (6'h1 == _T_198) begin
                                                          mem_1 <= _GEN_9;
                                                        end else begin
                                                          if (6'h1 == _T_193) begin
                                                            mem_1 <= _GEN_8;
                                                          end else begin
                                                            if (6'h1 == _T_188) begin
                                                              mem_1 <= _GEN_7;
                                                            end else begin
                                                              if (6'h1 == _T_183) begin
                                                                mem_1 <= _GEN_6;
                                                              end else begin
                                                                if (6'h1 == _T_178) begin
                                                                  mem_1 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h1 == _T_173) begin
                                                                    mem_1 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h1 == _T_168) begin
                                                                      mem_1 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h1 == _T_163) begin
                                                                        mem_1 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h1 == _T_158) begin
                                                                          mem_1 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h1 == _T_153) begin
                                                                            mem_1 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h1 == _T_308) begin
            mem_1 <= _GEN_31;
          end else begin
            if (6'h1 == _T_303) begin
              mem_1 <= _GEN_30;
            end else begin
              if (6'h1 == _T_298) begin
                mem_1 <= _GEN_29;
              end else begin
                if (6'h1 == _T_293) begin
                  mem_1 <= _GEN_28;
                end else begin
                  if (6'h1 == _T_288) begin
                    mem_1 <= _GEN_27;
                  end else begin
                    if (6'h1 == _T_283) begin
                      mem_1 <= _GEN_26;
                    end else begin
                      if (6'h1 == _T_278) begin
                        mem_1 <= _GEN_25;
                      end else begin
                        if (6'h1 == _T_273) begin
                          mem_1 <= _GEN_24;
                        end else begin
                          if (6'h1 == _T_268) begin
                            mem_1 <= _GEN_23;
                          end else begin
                            if (6'h1 == _T_263) begin
                              mem_1 <= _GEN_22;
                            end else begin
                              if (6'h1 == _T_258) begin
                                mem_1 <= _GEN_21;
                              end else begin
                                if (6'h1 == _T_253) begin
                                  mem_1 <= _GEN_20;
                                end else begin
                                  if (6'h1 == _T_248) begin
                                    mem_1 <= _GEN_19;
                                  end else begin
                                    if (6'h1 == _T_243) begin
                                      mem_1 <= _GEN_18;
                                    end else begin
                                      if (6'h1 == _T_238) begin
                                        mem_1 <= _GEN_17;
                                      end else begin
                                        if (6'h1 == _T_233) begin
                                          mem_1 <= _GEN_16;
                                        end else begin
                                          if (6'h1 == _T_228) begin
                                            mem_1 <= _GEN_15;
                                          end else begin
                                            if (6'h1 == _T_223) begin
                                              mem_1 <= _GEN_14;
                                            end else begin
                                              if (6'h1 == _T_218) begin
                                                mem_1 <= _GEN_13;
                                              end else begin
                                                if (6'h1 == _T_213) begin
                                                  mem_1 <= _GEN_12;
                                                end else begin
                                                  if (6'h1 == _T_208) begin
                                                    mem_1 <= _GEN_11;
                                                  end else begin
                                                    if (6'h1 == _T_203) begin
                                                      mem_1 <= _GEN_10;
                                                    end else begin
                                                      if (6'h1 == _T_198) begin
                                                        mem_1 <= _GEN_9;
                                                      end else begin
                                                        if (6'h1 == _T_193) begin
                                                          mem_1 <= _GEN_8;
                                                        end else begin
                                                          if (6'h1 == _T_188) begin
                                                            mem_1 <= _GEN_7;
                                                          end else begin
                                                            if (6'h1 == _T_183) begin
                                                              mem_1 <= _GEN_6;
                                                            end else begin
                                                              if (6'h1 == _T_178) begin
                                                                mem_1 <= _GEN_5;
                                                              end else begin
                                                                if (6'h1 == _T_173) begin
                                                                  mem_1 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h1 == _T_168) begin
                                                                    mem_1 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h1 == _T_163) begin
                                                                      mem_1 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h1 == _T_158) begin
                                                                        mem_1 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h1 == _T_153) begin
                                                                          mem_1 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h1 == _T_308) begin
          mem_1 <= _GEN_31;
        end else begin
          if (6'h1 == _T_303) begin
            mem_1 <= _GEN_30;
          end else begin
            if (6'h1 == _T_298) begin
              mem_1 <= _GEN_29;
            end else begin
              if (6'h1 == _T_293) begin
                mem_1 <= _GEN_28;
              end else begin
                if (6'h1 == _T_288) begin
                  mem_1 <= _GEN_27;
                end else begin
                  if (6'h1 == _T_283) begin
                    mem_1 <= _GEN_26;
                  end else begin
                    if (6'h1 == _T_278) begin
                      mem_1 <= _GEN_25;
                    end else begin
                      if (6'h1 == _T_273) begin
                        mem_1 <= _GEN_24;
                      end else begin
                        if (6'h1 == _T_268) begin
                          mem_1 <= _GEN_23;
                        end else begin
                          if (6'h1 == _T_263) begin
                            mem_1 <= _GEN_22;
                          end else begin
                            if (6'h1 == _T_258) begin
                              mem_1 <= _GEN_21;
                            end else begin
                              if (6'h1 == _T_253) begin
                                mem_1 <= _GEN_20;
                              end else begin
                                if (6'h1 == _T_248) begin
                                  mem_1 <= _GEN_19;
                                end else begin
                                  if (6'h1 == _T_243) begin
                                    mem_1 <= _GEN_18;
                                  end else begin
                                    if (6'h1 == _T_238) begin
                                      mem_1 <= _GEN_17;
                                    end else begin
                                      if (6'h1 == _T_233) begin
                                        mem_1 <= _GEN_16;
                                      end else begin
                                        if (6'h1 == _T_228) begin
                                          mem_1 <= _GEN_15;
                                        end else begin
                                          if (6'h1 == _T_223) begin
                                            mem_1 <= _GEN_14;
                                          end else begin
                                            if (6'h1 == _T_218) begin
                                              mem_1 <= _GEN_13;
                                            end else begin
                                              if (6'h1 == _T_213) begin
                                                mem_1 <= _GEN_12;
                                              end else begin
                                                if (6'h1 == _T_208) begin
                                                  mem_1 <= _GEN_11;
                                                end else begin
                                                  if (6'h1 == _T_203) begin
                                                    mem_1 <= _GEN_10;
                                                  end else begin
                                                    if (6'h1 == _T_198) begin
                                                      mem_1 <= _GEN_9;
                                                    end else begin
                                                      if (6'h1 == _T_193) begin
                                                        mem_1 <= _GEN_8;
                                                      end else begin
                                                        if (6'h1 == _T_188) begin
                                                          mem_1 <= _GEN_7;
                                                        end else begin
                                                          if (6'h1 == _T_183) begin
                                                            mem_1 <= _GEN_6;
                                                          end else begin
                                                            if (6'h1 == _T_178) begin
                                                              mem_1 <= _GEN_5;
                                                            end else begin
                                                              if (6'h1 == _T_173) begin
                                                                mem_1 <= _GEN_4;
                                                              end else begin
                                                                if (6'h1 == _T_168) begin
                                                                  mem_1 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h1 == _T_163) begin
                                                                    mem_1 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h1 == _T_158) begin
                                                                      mem_1 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h1 == _T_153) begin
                                                                        mem_1 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h2 == wPos) begin
            mem_2 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h2 == _T_308) begin
                mem_2 <= _GEN_31;
              end else begin
                if (6'h2 == _T_303) begin
                  mem_2 <= _GEN_30;
                end else begin
                  if (6'h2 == _T_298) begin
                    mem_2 <= _GEN_29;
                  end else begin
                    if (6'h2 == _T_293) begin
                      mem_2 <= _GEN_28;
                    end else begin
                      if (6'h2 == _T_288) begin
                        mem_2 <= _GEN_27;
                      end else begin
                        if (6'h2 == _T_283) begin
                          mem_2 <= _GEN_26;
                        end else begin
                          if (6'h2 == _T_278) begin
                            mem_2 <= _GEN_25;
                          end else begin
                            if (6'h2 == _T_273) begin
                              mem_2 <= _GEN_24;
                            end else begin
                              if (6'h2 == _T_268) begin
                                mem_2 <= _GEN_23;
                              end else begin
                                if (6'h2 == _T_263) begin
                                  mem_2 <= _GEN_22;
                                end else begin
                                  if (6'h2 == _T_258) begin
                                    mem_2 <= _GEN_21;
                                  end else begin
                                    if (6'h2 == _T_253) begin
                                      mem_2 <= _GEN_20;
                                    end else begin
                                      if (6'h2 == _T_248) begin
                                        mem_2 <= _GEN_19;
                                      end else begin
                                        if (6'h2 == _T_243) begin
                                          mem_2 <= _GEN_18;
                                        end else begin
                                          if (6'h2 == _T_238) begin
                                            mem_2 <= _GEN_17;
                                          end else begin
                                            if (6'h2 == _T_233) begin
                                              mem_2 <= _GEN_16;
                                            end else begin
                                              if (6'h2 == _T_228) begin
                                                mem_2 <= _GEN_15;
                                              end else begin
                                                if (6'h2 == _T_223) begin
                                                  mem_2 <= _GEN_14;
                                                end else begin
                                                  if (6'h2 == _T_218) begin
                                                    mem_2 <= _GEN_13;
                                                  end else begin
                                                    if (6'h2 == _T_213) begin
                                                      mem_2 <= _GEN_12;
                                                    end else begin
                                                      if (6'h2 == _T_208) begin
                                                        mem_2 <= _GEN_11;
                                                      end else begin
                                                        if (6'h2 == _T_203) begin
                                                          mem_2 <= _GEN_10;
                                                        end else begin
                                                          if (6'h2 == _T_198) begin
                                                            mem_2 <= _GEN_9;
                                                          end else begin
                                                            if (6'h2 == _T_193) begin
                                                              mem_2 <= _GEN_8;
                                                            end else begin
                                                              if (6'h2 == _T_188) begin
                                                                mem_2 <= _GEN_7;
                                                              end else begin
                                                                if (6'h2 == _T_183) begin
                                                                  mem_2 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h2 == _T_178) begin
                                                                    mem_2 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h2 == _T_173) begin
                                                                      mem_2 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h2 == _T_168) begin
                                                                        mem_2 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h2 == _T_163) begin
                                                                          mem_2 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h2 == _T_158) begin
                                                                            mem_2 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h2 == _T_153) begin
                                                                              mem_2 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h2 == _T_308) begin
              mem_2 <= _GEN_31;
            end else begin
              if (6'h2 == _T_303) begin
                mem_2 <= _GEN_30;
              end else begin
                if (6'h2 == _T_298) begin
                  mem_2 <= _GEN_29;
                end else begin
                  if (6'h2 == _T_293) begin
                    mem_2 <= _GEN_28;
                  end else begin
                    if (6'h2 == _T_288) begin
                      mem_2 <= _GEN_27;
                    end else begin
                      if (6'h2 == _T_283) begin
                        mem_2 <= _GEN_26;
                      end else begin
                        if (6'h2 == _T_278) begin
                          mem_2 <= _GEN_25;
                        end else begin
                          if (6'h2 == _T_273) begin
                            mem_2 <= _GEN_24;
                          end else begin
                            if (6'h2 == _T_268) begin
                              mem_2 <= _GEN_23;
                            end else begin
                              if (6'h2 == _T_263) begin
                                mem_2 <= _GEN_22;
                              end else begin
                                if (6'h2 == _T_258) begin
                                  mem_2 <= _GEN_21;
                                end else begin
                                  if (6'h2 == _T_253) begin
                                    mem_2 <= _GEN_20;
                                  end else begin
                                    if (6'h2 == _T_248) begin
                                      mem_2 <= _GEN_19;
                                    end else begin
                                      if (6'h2 == _T_243) begin
                                        mem_2 <= _GEN_18;
                                      end else begin
                                        if (6'h2 == _T_238) begin
                                          mem_2 <= _GEN_17;
                                        end else begin
                                          if (6'h2 == _T_233) begin
                                            mem_2 <= _GEN_16;
                                          end else begin
                                            if (6'h2 == _T_228) begin
                                              mem_2 <= _GEN_15;
                                            end else begin
                                              if (6'h2 == _T_223) begin
                                                mem_2 <= _GEN_14;
                                              end else begin
                                                if (6'h2 == _T_218) begin
                                                  mem_2 <= _GEN_13;
                                                end else begin
                                                  if (6'h2 == _T_213) begin
                                                    mem_2 <= _GEN_12;
                                                  end else begin
                                                    if (6'h2 == _T_208) begin
                                                      mem_2 <= _GEN_11;
                                                    end else begin
                                                      if (6'h2 == _T_203) begin
                                                        mem_2 <= _GEN_10;
                                                      end else begin
                                                        if (6'h2 == _T_198) begin
                                                          mem_2 <= _GEN_9;
                                                        end else begin
                                                          if (6'h2 == _T_193) begin
                                                            mem_2 <= _GEN_8;
                                                          end else begin
                                                            if (6'h2 == _T_188) begin
                                                              mem_2 <= _GEN_7;
                                                            end else begin
                                                              if (6'h2 == _T_183) begin
                                                                mem_2 <= _GEN_6;
                                                              end else begin
                                                                if (6'h2 == _T_178) begin
                                                                  mem_2 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h2 == _T_173) begin
                                                                    mem_2 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h2 == _T_168) begin
                                                                      mem_2 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h2 == _T_163) begin
                                                                        mem_2 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h2 == _T_158) begin
                                                                          mem_2 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h2 == _T_153) begin
                                                                            mem_2 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h2 == _T_308) begin
            mem_2 <= _GEN_31;
          end else begin
            if (6'h2 == _T_303) begin
              mem_2 <= _GEN_30;
            end else begin
              if (6'h2 == _T_298) begin
                mem_2 <= _GEN_29;
              end else begin
                if (6'h2 == _T_293) begin
                  mem_2 <= _GEN_28;
                end else begin
                  if (6'h2 == _T_288) begin
                    mem_2 <= _GEN_27;
                  end else begin
                    if (6'h2 == _T_283) begin
                      mem_2 <= _GEN_26;
                    end else begin
                      if (6'h2 == _T_278) begin
                        mem_2 <= _GEN_25;
                      end else begin
                        if (6'h2 == _T_273) begin
                          mem_2 <= _GEN_24;
                        end else begin
                          if (6'h2 == _T_268) begin
                            mem_2 <= _GEN_23;
                          end else begin
                            if (6'h2 == _T_263) begin
                              mem_2 <= _GEN_22;
                            end else begin
                              if (6'h2 == _T_258) begin
                                mem_2 <= _GEN_21;
                              end else begin
                                if (6'h2 == _T_253) begin
                                  mem_2 <= _GEN_20;
                                end else begin
                                  if (6'h2 == _T_248) begin
                                    mem_2 <= _GEN_19;
                                  end else begin
                                    if (6'h2 == _T_243) begin
                                      mem_2 <= _GEN_18;
                                    end else begin
                                      if (6'h2 == _T_238) begin
                                        mem_2 <= _GEN_17;
                                      end else begin
                                        if (6'h2 == _T_233) begin
                                          mem_2 <= _GEN_16;
                                        end else begin
                                          if (6'h2 == _T_228) begin
                                            mem_2 <= _GEN_15;
                                          end else begin
                                            if (6'h2 == _T_223) begin
                                              mem_2 <= _GEN_14;
                                            end else begin
                                              if (6'h2 == _T_218) begin
                                                mem_2 <= _GEN_13;
                                              end else begin
                                                if (6'h2 == _T_213) begin
                                                  mem_2 <= _GEN_12;
                                                end else begin
                                                  if (6'h2 == _T_208) begin
                                                    mem_2 <= _GEN_11;
                                                  end else begin
                                                    if (6'h2 == _T_203) begin
                                                      mem_2 <= _GEN_10;
                                                    end else begin
                                                      if (6'h2 == _T_198) begin
                                                        mem_2 <= _GEN_9;
                                                      end else begin
                                                        if (6'h2 == _T_193) begin
                                                          mem_2 <= _GEN_8;
                                                        end else begin
                                                          if (6'h2 == _T_188) begin
                                                            mem_2 <= _GEN_7;
                                                          end else begin
                                                            if (6'h2 == _T_183) begin
                                                              mem_2 <= _GEN_6;
                                                            end else begin
                                                              if (6'h2 == _T_178) begin
                                                                mem_2 <= _GEN_5;
                                                              end else begin
                                                                if (6'h2 == _T_173) begin
                                                                  mem_2 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h2 == _T_168) begin
                                                                    mem_2 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h2 == _T_163) begin
                                                                      mem_2 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h2 == _T_158) begin
                                                                        mem_2 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h2 == _T_153) begin
                                                                          mem_2 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h2 == _T_308) begin
          mem_2 <= _GEN_31;
        end else begin
          if (6'h2 == _T_303) begin
            mem_2 <= _GEN_30;
          end else begin
            if (6'h2 == _T_298) begin
              mem_2 <= _GEN_29;
            end else begin
              if (6'h2 == _T_293) begin
                mem_2 <= _GEN_28;
              end else begin
                if (6'h2 == _T_288) begin
                  mem_2 <= _GEN_27;
                end else begin
                  if (6'h2 == _T_283) begin
                    mem_2 <= _GEN_26;
                  end else begin
                    if (6'h2 == _T_278) begin
                      mem_2 <= _GEN_25;
                    end else begin
                      if (6'h2 == _T_273) begin
                        mem_2 <= _GEN_24;
                      end else begin
                        if (6'h2 == _T_268) begin
                          mem_2 <= _GEN_23;
                        end else begin
                          if (6'h2 == _T_263) begin
                            mem_2 <= _GEN_22;
                          end else begin
                            if (6'h2 == _T_258) begin
                              mem_2 <= _GEN_21;
                            end else begin
                              if (6'h2 == _T_253) begin
                                mem_2 <= _GEN_20;
                              end else begin
                                if (6'h2 == _T_248) begin
                                  mem_2 <= _GEN_19;
                                end else begin
                                  if (6'h2 == _T_243) begin
                                    mem_2 <= _GEN_18;
                                  end else begin
                                    if (6'h2 == _T_238) begin
                                      mem_2 <= _GEN_17;
                                    end else begin
                                      if (6'h2 == _T_233) begin
                                        mem_2 <= _GEN_16;
                                      end else begin
                                        if (6'h2 == _T_228) begin
                                          mem_2 <= _GEN_15;
                                        end else begin
                                          if (6'h2 == _T_223) begin
                                            mem_2 <= _GEN_14;
                                          end else begin
                                            if (6'h2 == _T_218) begin
                                              mem_2 <= _GEN_13;
                                            end else begin
                                              if (6'h2 == _T_213) begin
                                                mem_2 <= _GEN_12;
                                              end else begin
                                                if (6'h2 == _T_208) begin
                                                  mem_2 <= _GEN_11;
                                                end else begin
                                                  if (6'h2 == _T_203) begin
                                                    mem_2 <= _GEN_10;
                                                  end else begin
                                                    if (6'h2 == _T_198) begin
                                                      mem_2 <= _GEN_9;
                                                    end else begin
                                                      if (6'h2 == _T_193) begin
                                                        mem_2 <= _GEN_8;
                                                      end else begin
                                                        if (6'h2 == _T_188) begin
                                                          mem_2 <= _GEN_7;
                                                        end else begin
                                                          if (6'h2 == _T_183) begin
                                                            mem_2 <= _GEN_6;
                                                          end else begin
                                                            if (6'h2 == _T_178) begin
                                                              mem_2 <= _GEN_5;
                                                            end else begin
                                                              if (6'h2 == _T_173) begin
                                                                mem_2 <= _GEN_4;
                                                              end else begin
                                                                if (6'h2 == _T_168) begin
                                                                  mem_2 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h2 == _T_163) begin
                                                                    mem_2 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h2 == _T_158) begin
                                                                      mem_2 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h2 == _T_153) begin
                                                                        mem_2 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h3 == wPos) begin
            mem_3 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h3 == _T_308) begin
                mem_3 <= _GEN_31;
              end else begin
                if (6'h3 == _T_303) begin
                  mem_3 <= _GEN_30;
                end else begin
                  if (6'h3 == _T_298) begin
                    mem_3 <= _GEN_29;
                  end else begin
                    if (6'h3 == _T_293) begin
                      mem_3 <= _GEN_28;
                    end else begin
                      if (6'h3 == _T_288) begin
                        mem_3 <= _GEN_27;
                      end else begin
                        if (6'h3 == _T_283) begin
                          mem_3 <= _GEN_26;
                        end else begin
                          if (6'h3 == _T_278) begin
                            mem_3 <= _GEN_25;
                          end else begin
                            if (6'h3 == _T_273) begin
                              mem_3 <= _GEN_24;
                            end else begin
                              if (6'h3 == _T_268) begin
                                mem_3 <= _GEN_23;
                              end else begin
                                if (6'h3 == _T_263) begin
                                  mem_3 <= _GEN_22;
                                end else begin
                                  if (6'h3 == _T_258) begin
                                    mem_3 <= _GEN_21;
                                  end else begin
                                    if (6'h3 == _T_253) begin
                                      mem_3 <= _GEN_20;
                                    end else begin
                                      if (6'h3 == _T_248) begin
                                        mem_3 <= _GEN_19;
                                      end else begin
                                        if (6'h3 == _T_243) begin
                                          mem_3 <= _GEN_18;
                                        end else begin
                                          if (6'h3 == _T_238) begin
                                            mem_3 <= _GEN_17;
                                          end else begin
                                            if (6'h3 == _T_233) begin
                                              mem_3 <= _GEN_16;
                                            end else begin
                                              if (6'h3 == _T_228) begin
                                                mem_3 <= _GEN_15;
                                              end else begin
                                                if (6'h3 == _T_223) begin
                                                  mem_3 <= _GEN_14;
                                                end else begin
                                                  if (6'h3 == _T_218) begin
                                                    mem_3 <= _GEN_13;
                                                  end else begin
                                                    if (6'h3 == _T_213) begin
                                                      mem_3 <= _GEN_12;
                                                    end else begin
                                                      if (6'h3 == _T_208) begin
                                                        mem_3 <= _GEN_11;
                                                      end else begin
                                                        if (6'h3 == _T_203) begin
                                                          mem_3 <= _GEN_10;
                                                        end else begin
                                                          if (6'h3 == _T_198) begin
                                                            mem_3 <= _GEN_9;
                                                          end else begin
                                                            if (6'h3 == _T_193) begin
                                                              mem_3 <= _GEN_8;
                                                            end else begin
                                                              if (6'h3 == _T_188) begin
                                                                mem_3 <= _GEN_7;
                                                              end else begin
                                                                if (6'h3 == _T_183) begin
                                                                  mem_3 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h3 == _T_178) begin
                                                                    mem_3 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h3 == _T_173) begin
                                                                      mem_3 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h3 == _T_168) begin
                                                                        mem_3 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h3 == _T_163) begin
                                                                          mem_3 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h3 == _T_158) begin
                                                                            mem_3 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h3 == _T_153) begin
                                                                              mem_3 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h3 == _T_308) begin
              mem_3 <= _GEN_31;
            end else begin
              if (6'h3 == _T_303) begin
                mem_3 <= _GEN_30;
              end else begin
                if (6'h3 == _T_298) begin
                  mem_3 <= _GEN_29;
                end else begin
                  if (6'h3 == _T_293) begin
                    mem_3 <= _GEN_28;
                  end else begin
                    if (6'h3 == _T_288) begin
                      mem_3 <= _GEN_27;
                    end else begin
                      if (6'h3 == _T_283) begin
                        mem_3 <= _GEN_26;
                      end else begin
                        if (6'h3 == _T_278) begin
                          mem_3 <= _GEN_25;
                        end else begin
                          if (6'h3 == _T_273) begin
                            mem_3 <= _GEN_24;
                          end else begin
                            if (6'h3 == _T_268) begin
                              mem_3 <= _GEN_23;
                            end else begin
                              if (6'h3 == _T_263) begin
                                mem_3 <= _GEN_22;
                              end else begin
                                if (6'h3 == _T_258) begin
                                  mem_3 <= _GEN_21;
                                end else begin
                                  if (6'h3 == _T_253) begin
                                    mem_3 <= _GEN_20;
                                  end else begin
                                    if (6'h3 == _T_248) begin
                                      mem_3 <= _GEN_19;
                                    end else begin
                                      if (6'h3 == _T_243) begin
                                        mem_3 <= _GEN_18;
                                      end else begin
                                        if (6'h3 == _T_238) begin
                                          mem_3 <= _GEN_17;
                                        end else begin
                                          if (6'h3 == _T_233) begin
                                            mem_3 <= _GEN_16;
                                          end else begin
                                            if (6'h3 == _T_228) begin
                                              mem_3 <= _GEN_15;
                                            end else begin
                                              if (6'h3 == _T_223) begin
                                                mem_3 <= _GEN_14;
                                              end else begin
                                                if (6'h3 == _T_218) begin
                                                  mem_3 <= _GEN_13;
                                                end else begin
                                                  if (6'h3 == _T_213) begin
                                                    mem_3 <= _GEN_12;
                                                  end else begin
                                                    if (6'h3 == _T_208) begin
                                                      mem_3 <= _GEN_11;
                                                    end else begin
                                                      if (6'h3 == _T_203) begin
                                                        mem_3 <= _GEN_10;
                                                      end else begin
                                                        if (6'h3 == _T_198) begin
                                                          mem_3 <= _GEN_9;
                                                        end else begin
                                                          if (6'h3 == _T_193) begin
                                                            mem_3 <= _GEN_8;
                                                          end else begin
                                                            if (6'h3 == _T_188) begin
                                                              mem_3 <= _GEN_7;
                                                            end else begin
                                                              if (6'h3 == _T_183) begin
                                                                mem_3 <= _GEN_6;
                                                              end else begin
                                                                if (6'h3 == _T_178) begin
                                                                  mem_3 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h3 == _T_173) begin
                                                                    mem_3 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h3 == _T_168) begin
                                                                      mem_3 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h3 == _T_163) begin
                                                                        mem_3 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h3 == _T_158) begin
                                                                          mem_3 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h3 == _T_153) begin
                                                                            mem_3 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h3 == _T_308) begin
            mem_3 <= _GEN_31;
          end else begin
            if (6'h3 == _T_303) begin
              mem_3 <= _GEN_30;
            end else begin
              if (6'h3 == _T_298) begin
                mem_3 <= _GEN_29;
              end else begin
                if (6'h3 == _T_293) begin
                  mem_3 <= _GEN_28;
                end else begin
                  if (6'h3 == _T_288) begin
                    mem_3 <= _GEN_27;
                  end else begin
                    if (6'h3 == _T_283) begin
                      mem_3 <= _GEN_26;
                    end else begin
                      if (6'h3 == _T_278) begin
                        mem_3 <= _GEN_25;
                      end else begin
                        if (6'h3 == _T_273) begin
                          mem_3 <= _GEN_24;
                        end else begin
                          if (6'h3 == _T_268) begin
                            mem_3 <= _GEN_23;
                          end else begin
                            if (6'h3 == _T_263) begin
                              mem_3 <= _GEN_22;
                            end else begin
                              if (6'h3 == _T_258) begin
                                mem_3 <= _GEN_21;
                              end else begin
                                if (6'h3 == _T_253) begin
                                  mem_3 <= _GEN_20;
                                end else begin
                                  if (6'h3 == _T_248) begin
                                    mem_3 <= _GEN_19;
                                  end else begin
                                    if (6'h3 == _T_243) begin
                                      mem_3 <= _GEN_18;
                                    end else begin
                                      if (6'h3 == _T_238) begin
                                        mem_3 <= _GEN_17;
                                      end else begin
                                        if (6'h3 == _T_233) begin
                                          mem_3 <= _GEN_16;
                                        end else begin
                                          if (6'h3 == _T_228) begin
                                            mem_3 <= _GEN_15;
                                          end else begin
                                            if (6'h3 == _T_223) begin
                                              mem_3 <= _GEN_14;
                                            end else begin
                                              if (6'h3 == _T_218) begin
                                                mem_3 <= _GEN_13;
                                              end else begin
                                                if (6'h3 == _T_213) begin
                                                  mem_3 <= _GEN_12;
                                                end else begin
                                                  if (6'h3 == _T_208) begin
                                                    mem_3 <= _GEN_11;
                                                  end else begin
                                                    if (6'h3 == _T_203) begin
                                                      mem_3 <= _GEN_10;
                                                    end else begin
                                                      if (6'h3 == _T_198) begin
                                                        mem_3 <= _GEN_9;
                                                      end else begin
                                                        if (6'h3 == _T_193) begin
                                                          mem_3 <= _GEN_8;
                                                        end else begin
                                                          if (6'h3 == _T_188) begin
                                                            mem_3 <= _GEN_7;
                                                          end else begin
                                                            if (6'h3 == _T_183) begin
                                                              mem_3 <= _GEN_6;
                                                            end else begin
                                                              if (6'h3 == _T_178) begin
                                                                mem_3 <= _GEN_5;
                                                              end else begin
                                                                if (6'h3 == _T_173) begin
                                                                  mem_3 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h3 == _T_168) begin
                                                                    mem_3 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h3 == _T_163) begin
                                                                      mem_3 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h3 == _T_158) begin
                                                                        mem_3 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h3 == _T_153) begin
                                                                          mem_3 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h3 == _T_308) begin
          mem_3 <= _GEN_31;
        end else begin
          if (6'h3 == _T_303) begin
            mem_3 <= _GEN_30;
          end else begin
            if (6'h3 == _T_298) begin
              mem_3 <= _GEN_29;
            end else begin
              if (6'h3 == _T_293) begin
                mem_3 <= _GEN_28;
              end else begin
                if (6'h3 == _T_288) begin
                  mem_3 <= _GEN_27;
                end else begin
                  if (6'h3 == _T_283) begin
                    mem_3 <= _GEN_26;
                  end else begin
                    if (6'h3 == _T_278) begin
                      mem_3 <= _GEN_25;
                    end else begin
                      if (6'h3 == _T_273) begin
                        mem_3 <= _GEN_24;
                      end else begin
                        if (6'h3 == _T_268) begin
                          mem_3 <= _GEN_23;
                        end else begin
                          if (6'h3 == _T_263) begin
                            mem_3 <= _GEN_22;
                          end else begin
                            if (6'h3 == _T_258) begin
                              mem_3 <= _GEN_21;
                            end else begin
                              if (6'h3 == _T_253) begin
                                mem_3 <= _GEN_20;
                              end else begin
                                if (6'h3 == _T_248) begin
                                  mem_3 <= _GEN_19;
                                end else begin
                                  if (6'h3 == _T_243) begin
                                    mem_3 <= _GEN_18;
                                  end else begin
                                    if (6'h3 == _T_238) begin
                                      mem_3 <= _GEN_17;
                                    end else begin
                                      if (6'h3 == _T_233) begin
                                        mem_3 <= _GEN_16;
                                      end else begin
                                        if (6'h3 == _T_228) begin
                                          mem_3 <= _GEN_15;
                                        end else begin
                                          if (6'h3 == _T_223) begin
                                            mem_3 <= _GEN_14;
                                          end else begin
                                            if (6'h3 == _T_218) begin
                                              mem_3 <= _GEN_13;
                                            end else begin
                                              if (6'h3 == _T_213) begin
                                                mem_3 <= _GEN_12;
                                              end else begin
                                                if (6'h3 == _T_208) begin
                                                  mem_3 <= _GEN_11;
                                                end else begin
                                                  if (6'h3 == _T_203) begin
                                                    mem_3 <= _GEN_10;
                                                  end else begin
                                                    if (6'h3 == _T_198) begin
                                                      mem_3 <= _GEN_9;
                                                    end else begin
                                                      if (6'h3 == _T_193) begin
                                                        mem_3 <= _GEN_8;
                                                      end else begin
                                                        if (6'h3 == _T_188) begin
                                                          mem_3 <= _GEN_7;
                                                        end else begin
                                                          if (6'h3 == _T_183) begin
                                                            mem_3 <= _GEN_6;
                                                          end else begin
                                                            if (6'h3 == _T_178) begin
                                                              mem_3 <= _GEN_5;
                                                            end else begin
                                                              if (6'h3 == _T_173) begin
                                                                mem_3 <= _GEN_4;
                                                              end else begin
                                                                if (6'h3 == _T_168) begin
                                                                  mem_3 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h3 == _T_163) begin
                                                                    mem_3 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h3 == _T_158) begin
                                                                      mem_3 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h3 == _T_153) begin
                                                                        mem_3 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h4 == wPos) begin
            mem_4 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h4 == _T_308) begin
                mem_4 <= _GEN_31;
              end else begin
                if (6'h4 == _T_303) begin
                  mem_4 <= _GEN_30;
                end else begin
                  if (6'h4 == _T_298) begin
                    mem_4 <= _GEN_29;
                  end else begin
                    if (6'h4 == _T_293) begin
                      mem_4 <= _GEN_28;
                    end else begin
                      if (6'h4 == _T_288) begin
                        mem_4 <= _GEN_27;
                      end else begin
                        if (6'h4 == _T_283) begin
                          mem_4 <= _GEN_26;
                        end else begin
                          if (6'h4 == _T_278) begin
                            mem_4 <= _GEN_25;
                          end else begin
                            if (6'h4 == _T_273) begin
                              mem_4 <= _GEN_24;
                            end else begin
                              if (6'h4 == _T_268) begin
                                mem_4 <= _GEN_23;
                              end else begin
                                if (6'h4 == _T_263) begin
                                  mem_4 <= _GEN_22;
                                end else begin
                                  if (6'h4 == _T_258) begin
                                    mem_4 <= _GEN_21;
                                  end else begin
                                    if (6'h4 == _T_253) begin
                                      mem_4 <= _GEN_20;
                                    end else begin
                                      if (6'h4 == _T_248) begin
                                        mem_4 <= _GEN_19;
                                      end else begin
                                        if (6'h4 == _T_243) begin
                                          mem_4 <= _GEN_18;
                                        end else begin
                                          if (6'h4 == _T_238) begin
                                            mem_4 <= _GEN_17;
                                          end else begin
                                            if (6'h4 == _T_233) begin
                                              mem_4 <= _GEN_16;
                                            end else begin
                                              if (6'h4 == _T_228) begin
                                                mem_4 <= _GEN_15;
                                              end else begin
                                                if (6'h4 == _T_223) begin
                                                  mem_4 <= _GEN_14;
                                                end else begin
                                                  if (6'h4 == _T_218) begin
                                                    mem_4 <= _GEN_13;
                                                  end else begin
                                                    if (6'h4 == _T_213) begin
                                                      mem_4 <= _GEN_12;
                                                    end else begin
                                                      if (6'h4 == _T_208) begin
                                                        mem_4 <= _GEN_11;
                                                      end else begin
                                                        if (6'h4 == _T_203) begin
                                                          mem_4 <= _GEN_10;
                                                        end else begin
                                                          if (6'h4 == _T_198) begin
                                                            mem_4 <= _GEN_9;
                                                          end else begin
                                                            if (6'h4 == _T_193) begin
                                                              mem_4 <= _GEN_8;
                                                            end else begin
                                                              if (6'h4 == _T_188) begin
                                                                mem_4 <= _GEN_7;
                                                              end else begin
                                                                if (6'h4 == _T_183) begin
                                                                  mem_4 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h4 == _T_178) begin
                                                                    mem_4 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h4 == _T_173) begin
                                                                      mem_4 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h4 == _T_168) begin
                                                                        mem_4 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h4 == _T_163) begin
                                                                          mem_4 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h4 == _T_158) begin
                                                                            mem_4 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h4 == _T_153) begin
                                                                              mem_4 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h4 == _T_308) begin
              mem_4 <= _GEN_31;
            end else begin
              if (6'h4 == _T_303) begin
                mem_4 <= _GEN_30;
              end else begin
                if (6'h4 == _T_298) begin
                  mem_4 <= _GEN_29;
                end else begin
                  if (6'h4 == _T_293) begin
                    mem_4 <= _GEN_28;
                  end else begin
                    if (6'h4 == _T_288) begin
                      mem_4 <= _GEN_27;
                    end else begin
                      if (6'h4 == _T_283) begin
                        mem_4 <= _GEN_26;
                      end else begin
                        if (6'h4 == _T_278) begin
                          mem_4 <= _GEN_25;
                        end else begin
                          if (6'h4 == _T_273) begin
                            mem_4 <= _GEN_24;
                          end else begin
                            if (6'h4 == _T_268) begin
                              mem_4 <= _GEN_23;
                            end else begin
                              if (6'h4 == _T_263) begin
                                mem_4 <= _GEN_22;
                              end else begin
                                if (6'h4 == _T_258) begin
                                  mem_4 <= _GEN_21;
                                end else begin
                                  if (6'h4 == _T_253) begin
                                    mem_4 <= _GEN_20;
                                  end else begin
                                    if (6'h4 == _T_248) begin
                                      mem_4 <= _GEN_19;
                                    end else begin
                                      if (6'h4 == _T_243) begin
                                        mem_4 <= _GEN_18;
                                      end else begin
                                        if (6'h4 == _T_238) begin
                                          mem_4 <= _GEN_17;
                                        end else begin
                                          if (6'h4 == _T_233) begin
                                            mem_4 <= _GEN_16;
                                          end else begin
                                            if (6'h4 == _T_228) begin
                                              mem_4 <= _GEN_15;
                                            end else begin
                                              if (6'h4 == _T_223) begin
                                                mem_4 <= _GEN_14;
                                              end else begin
                                                if (6'h4 == _T_218) begin
                                                  mem_4 <= _GEN_13;
                                                end else begin
                                                  if (6'h4 == _T_213) begin
                                                    mem_4 <= _GEN_12;
                                                  end else begin
                                                    if (6'h4 == _T_208) begin
                                                      mem_4 <= _GEN_11;
                                                    end else begin
                                                      if (6'h4 == _T_203) begin
                                                        mem_4 <= _GEN_10;
                                                      end else begin
                                                        if (6'h4 == _T_198) begin
                                                          mem_4 <= _GEN_9;
                                                        end else begin
                                                          if (6'h4 == _T_193) begin
                                                            mem_4 <= _GEN_8;
                                                          end else begin
                                                            if (6'h4 == _T_188) begin
                                                              mem_4 <= _GEN_7;
                                                            end else begin
                                                              if (6'h4 == _T_183) begin
                                                                mem_4 <= _GEN_6;
                                                              end else begin
                                                                if (6'h4 == _T_178) begin
                                                                  mem_4 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h4 == _T_173) begin
                                                                    mem_4 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h4 == _T_168) begin
                                                                      mem_4 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h4 == _T_163) begin
                                                                        mem_4 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h4 == _T_158) begin
                                                                          mem_4 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h4 == _T_153) begin
                                                                            mem_4 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h4 == _T_308) begin
            mem_4 <= _GEN_31;
          end else begin
            if (6'h4 == _T_303) begin
              mem_4 <= _GEN_30;
            end else begin
              if (6'h4 == _T_298) begin
                mem_4 <= _GEN_29;
              end else begin
                if (6'h4 == _T_293) begin
                  mem_4 <= _GEN_28;
                end else begin
                  if (6'h4 == _T_288) begin
                    mem_4 <= _GEN_27;
                  end else begin
                    if (6'h4 == _T_283) begin
                      mem_4 <= _GEN_26;
                    end else begin
                      if (6'h4 == _T_278) begin
                        mem_4 <= _GEN_25;
                      end else begin
                        if (6'h4 == _T_273) begin
                          mem_4 <= _GEN_24;
                        end else begin
                          if (6'h4 == _T_268) begin
                            mem_4 <= _GEN_23;
                          end else begin
                            if (6'h4 == _T_263) begin
                              mem_4 <= _GEN_22;
                            end else begin
                              if (6'h4 == _T_258) begin
                                mem_4 <= _GEN_21;
                              end else begin
                                if (6'h4 == _T_253) begin
                                  mem_4 <= _GEN_20;
                                end else begin
                                  if (6'h4 == _T_248) begin
                                    mem_4 <= _GEN_19;
                                  end else begin
                                    if (6'h4 == _T_243) begin
                                      mem_4 <= _GEN_18;
                                    end else begin
                                      if (6'h4 == _T_238) begin
                                        mem_4 <= _GEN_17;
                                      end else begin
                                        if (6'h4 == _T_233) begin
                                          mem_4 <= _GEN_16;
                                        end else begin
                                          if (6'h4 == _T_228) begin
                                            mem_4 <= _GEN_15;
                                          end else begin
                                            if (6'h4 == _T_223) begin
                                              mem_4 <= _GEN_14;
                                            end else begin
                                              if (6'h4 == _T_218) begin
                                                mem_4 <= _GEN_13;
                                              end else begin
                                                if (6'h4 == _T_213) begin
                                                  mem_4 <= _GEN_12;
                                                end else begin
                                                  if (6'h4 == _T_208) begin
                                                    mem_4 <= _GEN_11;
                                                  end else begin
                                                    if (6'h4 == _T_203) begin
                                                      mem_4 <= _GEN_10;
                                                    end else begin
                                                      if (6'h4 == _T_198) begin
                                                        mem_4 <= _GEN_9;
                                                      end else begin
                                                        if (6'h4 == _T_193) begin
                                                          mem_4 <= _GEN_8;
                                                        end else begin
                                                          if (6'h4 == _T_188) begin
                                                            mem_4 <= _GEN_7;
                                                          end else begin
                                                            if (6'h4 == _T_183) begin
                                                              mem_4 <= _GEN_6;
                                                            end else begin
                                                              if (6'h4 == _T_178) begin
                                                                mem_4 <= _GEN_5;
                                                              end else begin
                                                                if (6'h4 == _T_173) begin
                                                                  mem_4 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h4 == _T_168) begin
                                                                    mem_4 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h4 == _T_163) begin
                                                                      mem_4 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h4 == _T_158) begin
                                                                        mem_4 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h4 == _T_153) begin
                                                                          mem_4 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h4 == _T_308) begin
          mem_4 <= _GEN_31;
        end else begin
          if (6'h4 == _T_303) begin
            mem_4 <= _GEN_30;
          end else begin
            if (6'h4 == _T_298) begin
              mem_4 <= _GEN_29;
            end else begin
              if (6'h4 == _T_293) begin
                mem_4 <= _GEN_28;
              end else begin
                if (6'h4 == _T_288) begin
                  mem_4 <= _GEN_27;
                end else begin
                  if (6'h4 == _T_283) begin
                    mem_4 <= _GEN_26;
                  end else begin
                    if (6'h4 == _T_278) begin
                      mem_4 <= _GEN_25;
                    end else begin
                      if (6'h4 == _T_273) begin
                        mem_4 <= _GEN_24;
                      end else begin
                        if (6'h4 == _T_268) begin
                          mem_4 <= _GEN_23;
                        end else begin
                          if (6'h4 == _T_263) begin
                            mem_4 <= _GEN_22;
                          end else begin
                            if (6'h4 == _T_258) begin
                              mem_4 <= _GEN_21;
                            end else begin
                              if (6'h4 == _T_253) begin
                                mem_4 <= _GEN_20;
                              end else begin
                                if (6'h4 == _T_248) begin
                                  mem_4 <= _GEN_19;
                                end else begin
                                  if (6'h4 == _T_243) begin
                                    mem_4 <= _GEN_18;
                                  end else begin
                                    if (6'h4 == _T_238) begin
                                      mem_4 <= _GEN_17;
                                    end else begin
                                      if (6'h4 == _T_233) begin
                                        mem_4 <= _GEN_16;
                                      end else begin
                                        if (6'h4 == _T_228) begin
                                          mem_4 <= _GEN_15;
                                        end else begin
                                          if (6'h4 == _T_223) begin
                                            mem_4 <= _GEN_14;
                                          end else begin
                                            if (6'h4 == _T_218) begin
                                              mem_4 <= _GEN_13;
                                            end else begin
                                              if (6'h4 == _T_213) begin
                                                mem_4 <= _GEN_12;
                                              end else begin
                                                if (6'h4 == _T_208) begin
                                                  mem_4 <= _GEN_11;
                                                end else begin
                                                  if (6'h4 == _T_203) begin
                                                    mem_4 <= _GEN_10;
                                                  end else begin
                                                    if (6'h4 == _T_198) begin
                                                      mem_4 <= _GEN_9;
                                                    end else begin
                                                      if (6'h4 == _T_193) begin
                                                        mem_4 <= _GEN_8;
                                                      end else begin
                                                        if (6'h4 == _T_188) begin
                                                          mem_4 <= _GEN_7;
                                                        end else begin
                                                          if (6'h4 == _T_183) begin
                                                            mem_4 <= _GEN_6;
                                                          end else begin
                                                            if (6'h4 == _T_178) begin
                                                              mem_4 <= _GEN_5;
                                                            end else begin
                                                              if (6'h4 == _T_173) begin
                                                                mem_4 <= _GEN_4;
                                                              end else begin
                                                                if (6'h4 == _T_168) begin
                                                                  mem_4 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h4 == _T_163) begin
                                                                    mem_4 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h4 == _T_158) begin
                                                                      mem_4 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h4 == _T_153) begin
                                                                        mem_4 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h5 == wPos) begin
            mem_5 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h5 == _T_308) begin
                mem_5 <= _GEN_31;
              end else begin
                if (6'h5 == _T_303) begin
                  mem_5 <= _GEN_30;
                end else begin
                  if (6'h5 == _T_298) begin
                    mem_5 <= _GEN_29;
                  end else begin
                    if (6'h5 == _T_293) begin
                      mem_5 <= _GEN_28;
                    end else begin
                      if (6'h5 == _T_288) begin
                        mem_5 <= _GEN_27;
                      end else begin
                        if (6'h5 == _T_283) begin
                          mem_5 <= _GEN_26;
                        end else begin
                          if (6'h5 == _T_278) begin
                            mem_5 <= _GEN_25;
                          end else begin
                            if (6'h5 == _T_273) begin
                              mem_5 <= _GEN_24;
                            end else begin
                              if (6'h5 == _T_268) begin
                                mem_5 <= _GEN_23;
                              end else begin
                                if (6'h5 == _T_263) begin
                                  mem_5 <= _GEN_22;
                                end else begin
                                  if (6'h5 == _T_258) begin
                                    mem_5 <= _GEN_21;
                                  end else begin
                                    if (6'h5 == _T_253) begin
                                      mem_5 <= _GEN_20;
                                    end else begin
                                      if (6'h5 == _T_248) begin
                                        mem_5 <= _GEN_19;
                                      end else begin
                                        if (6'h5 == _T_243) begin
                                          mem_5 <= _GEN_18;
                                        end else begin
                                          if (6'h5 == _T_238) begin
                                            mem_5 <= _GEN_17;
                                          end else begin
                                            if (6'h5 == _T_233) begin
                                              mem_5 <= _GEN_16;
                                            end else begin
                                              if (6'h5 == _T_228) begin
                                                mem_5 <= _GEN_15;
                                              end else begin
                                                if (6'h5 == _T_223) begin
                                                  mem_5 <= _GEN_14;
                                                end else begin
                                                  if (6'h5 == _T_218) begin
                                                    mem_5 <= _GEN_13;
                                                  end else begin
                                                    if (6'h5 == _T_213) begin
                                                      mem_5 <= _GEN_12;
                                                    end else begin
                                                      if (6'h5 == _T_208) begin
                                                        mem_5 <= _GEN_11;
                                                      end else begin
                                                        if (6'h5 == _T_203) begin
                                                          mem_5 <= _GEN_10;
                                                        end else begin
                                                          if (6'h5 == _T_198) begin
                                                            mem_5 <= _GEN_9;
                                                          end else begin
                                                            if (6'h5 == _T_193) begin
                                                              mem_5 <= _GEN_8;
                                                            end else begin
                                                              if (6'h5 == _T_188) begin
                                                                mem_5 <= _GEN_7;
                                                              end else begin
                                                                if (6'h5 == _T_183) begin
                                                                  mem_5 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h5 == _T_178) begin
                                                                    mem_5 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h5 == _T_173) begin
                                                                      mem_5 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h5 == _T_168) begin
                                                                        mem_5 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h5 == _T_163) begin
                                                                          mem_5 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h5 == _T_158) begin
                                                                            mem_5 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h5 == _T_153) begin
                                                                              mem_5 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h5 == _T_308) begin
              mem_5 <= _GEN_31;
            end else begin
              if (6'h5 == _T_303) begin
                mem_5 <= _GEN_30;
              end else begin
                if (6'h5 == _T_298) begin
                  mem_5 <= _GEN_29;
                end else begin
                  if (6'h5 == _T_293) begin
                    mem_5 <= _GEN_28;
                  end else begin
                    if (6'h5 == _T_288) begin
                      mem_5 <= _GEN_27;
                    end else begin
                      if (6'h5 == _T_283) begin
                        mem_5 <= _GEN_26;
                      end else begin
                        if (6'h5 == _T_278) begin
                          mem_5 <= _GEN_25;
                        end else begin
                          if (6'h5 == _T_273) begin
                            mem_5 <= _GEN_24;
                          end else begin
                            if (6'h5 == _T_268) begin
                              mem_5 <= _GEN_23;
                            end else begin
                              if (6'h5 == _T_263) begin
                                mem_5 <= _GEN_22;
                              end else begin
                                if (6'h5 == _T_258) begin
                                  mem_5 <= _GEN_21;
                                end else begin
                                  if (6'h5 == _T_253) begin
                                    mem_5 <= _GEN_20;
                                  end else begin
                                    if (6'h5 == _T_248) begin
                                      mem_5 <= _GEN_19;
                                    end else begin
                                      if (6'h5 == _T_243) begin
                                        mem_5 <= _GEN_18;
                                      end else begin
                                        if (6'h5 == _T_238) begin
                                          mem_5 <= _GEN_17;
                                        end else begin
                                          if (6'h5 == _T_233) begin
                                            mem_5 <= _GEN_16;
                                          end else begin
                                            if (6'h5 == _T_228) begin
                                              mem_5 <= _GEN_15;
                                            end else begin
                                              if (6'h5 == _T_223) begin
                                                mem_5 <= _GEN_14;
                                              end else begin
                                                if (6'h5 == _T_218) begin
                                                  mem_5 <= _GEN_13;
                                                end else begin
                                                  if (6'h5 == _T_213) begin
                                                    mem_5 <= _GEN_12;
                                                  end else begin
                                                    if (6'h5 == _T_208) begin
                                                      mem_5 <= _GEN_11;
                                                    end else begin
                                                      if (6'h5 == _T_203) begin
                                                        mem_5 <= _GEN_10;
                                                      end else begin
                                                        if (6'h5 == _T_198) begin
                                                          mem_5 <= _GEN_9;
                                                        end else begin
                                                          if (6'h5 == _T_193) begin
                                                            mem_5 <= _GEN_8;
                                                          end else begin
                                                            if (6'h5 == _T_188) begin
                                                              mem_5 <= _GEN_7;
                                                            end else begin
                                                              if (6'h5 == _T_183) begin
                                                                mem_5 <= _GEN_6;
                                                              end else begin
                                                                if (6'h5 == _T_178) begin
                                                                  mem_5 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h5 == _T_173) begin
                                                                    mem_5 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h5 == _T_168) begin
                                                                      mem_5 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h5 == _T_163) begin
                                                                        mem_5 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h5 == _T_158) begin
                                                                          mem_5 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h5 == _T_153) begin
                                                                            mem_5 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h5 == _T_308) begin
            mem_5 <= _GEN_31;
          end else begin
            if (6'h5 == _T_303) begin
              mem_5 <= _GEN_30;
            end else begin
              if (6'h5 == _T_298) begin
                mem_5 <= _GEN_29;
              end else begin
                if (6'h5 == _T_293) begin
                  mem_5 <= _GEN_28;
                end else begin
                  if (6'h5 == _T_288) begin
                    mem_5 <= _GEN_27;
                  end else begin
                    if (6'h5 == _T_283) begin
                      mem_5 <= _GEN_26;
                    end else begin
                      if (6'h5 == _T_278) begin
                        mem_5 <= _GEN_25;
                      end else begin
                        if (6'h5 == _T_273) begin
                          mem_5 <= _GEN_24;
                        end else begin
                          if (6'h5 == _T_268) begin
                            mem_5 <= _GEN_23;
                          end else begin
                            if (6'h5 == _T_263) begin
                              mem_5 <= _GEN_22;
                            end else begin
                              if (6'h5 == _T_258) begin
                                mem_5 <= _GEN_21;
                              end else begin
                                if (6'h5 == _T_253) begin
                                  mem_5 <= _GEN_20;
                                end else begin
                                  if (6'h5 == _T_248) begin
                                    mem_5 <= _GEN_19;
                                  end else begin
                                    if (6'h5 == _T_243) begin
                                      mem_5 <= _GEN_18;
                                    end else begin
                                      if (6'h5 == _T_238) begin
                                        mem_5 <= _GEN_17;
                                      end else begin
                                        if (6'h5 == _T_233) begin
                                          mem_5 <= _GEN_16;
                                        end else begin
                                          if (6'h5 == _T_228) begin
                                            mem_5 <= _GEN_15;
                                          end else begin
                                            if (6'h5 == _T_223) begin
                                              mem_5 <= _GEN_14;
                                            end else begin
                                              if (6'h5 == _T_218) begin
                                                mem_5 <= _GEN_13;
                                              end else begin
                                                if (6'h5 == _T_213) begin
                                                  mem_5 <= _GEN_12;
                                                end else begin
                                                  if (6'h5 == _T_208) begin
                                                    mem_5 <= _GEN_11;
                                                  end else begin
                                                    if (6'h5 == _T_203) begin
                                                      mem_5 <= _GEN_10;
                                                    end else begin
                                                      if (6'h5 == _T_198) begin
                                                        mem_5 <= _GEN_9;
                                                      end else begin
                                                        if (6'h5 == _T_193) begin
                                                          mem_5 <= _GEN_8;
                                                        end else begin
                                                          if (6'h5 == _T_188) begin
                                                            mem_5 <= _GEN_7;
                                                          end else begin
                                                            if (6'h5 == _T_183) begin
                                                              mem_5 <= _GEN_6;
                                                            end else begin
                                                              if (6'h5 == _T_178) begin
                                                                mem_5 <= _GEN_5;
                                                              end else begin
                                                                if (6'h5 == _T_173) begin
                                                                  mem_5 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h5 == _T_168) begin
                                                                    mem_5 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h5 == _T_163) begin
                                                                      mem_5 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h5 == _T_158) begin
                                                                        mem_5 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h5 == _T_153) begin
                                                                          mem_5 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h5 == _T_308) begin
          mem_5 <= _GEN_31;
        end else begin
          if (6'h5 == _T_303) begin
            mem_5 <= _GEN_30;
          end else begin
            if (6'h5 == _T_298) begin
              mem_5 <= _GEN_29;
            end else begin
              if (6'h5 == _T_293) begin
                mem_5 <= _GEN_28;
              end else begin
                if (6'h5 == _T_288) begin
                  mem_5 <= _GEN_27;
                end else begin
                  if (6'h5 == _T_283) begin
                    mem_5 <= _GEN_26;
                  end else begin
                    if (6'h5 == _T_278) begin
                      mem_5 <= _GEN_25;
                    end else begin
                      if (6'h5 == _T_273) begin
                        mem_5 <= _GEN_24;
                      end else begin
                        if (6'h5 == _T_268) begin
                          mem_5 <= _GEN_23;
                        end else begin
                          if (6'h5 == _T_263) begin
                            mem_5 <= _GEN_22;
                          end else begin
                            if (6'h5 == _T_258) begin
                              mem_5 <= _GEN_21;
                            end else begin
                              if (6'h5 == _T_253) begin
                                mem_5 <= _GEN_20;
                              end else begin
                                if (6'h5 == _T_248) begin
                                  mem_5 <= _GEN_19;
                                end else begin
                                  if (6'h5 == _T_243) begin
                                    mem_5 <= _GEN_18;
                                  end else begin
                                    if (6'h5 == _T_238) begin
                                      mem_5 <= _GEN_17;
                                    end else begin
                                      if (6'h5 == _T_233) begin
                                        mem_5 <= _GEN_16;
                                      end else begin
                                        if (6'h5 == _T_228) begin
                                          mem_5 <= _GEN_15;
                                        end else begin
                                          if (6'h5 == _T_223) begin
                                            mem_5 <= _GEN_14;
                                          end else begin
                                            if (6'h5 == _T_218) begin
                                              mem_5 <= _GEN_13;
                                            end else begin
                                              if (6'h5 == _T_213) begin
                                                mem_5 <= _GEN_12;
                                              end else begin
                                                if (6'h5 == _T_208) begin
                                                  mem_5 <= _GEN_11;
                                                end else begin
                                                  if (6'h5 == _T_203) begin
                                                    mem_5 <= _GEN_10;
                                                  end else begin
                                                    if (6'h5 == _T_198) begin
                                                      mem_5 <= _GEN_9;
                                                    end else begin
                                                      if (6'h5 == _T_193) begin
                                                        mem_5 <= _GEN_8;
                                                      end else begin
                                                        if (6'h5 == _T_188) begin
                                                          mem_5 <= _GEN_7;
                                                        end else begin
                                                          if (6'h5 == _T_183) begin
                                                            mem_5 <= _GEN_6;
                                                          end else begin
                                                            if (6'h5 == _T_178) begin
                                                              mem_5 <= _GEN_5;
                                                            end else begin
                                                              if (6'h5 == _T_173) begin
                                                                mem_5 <= _GEN_4;
                                                              end else begin
                                                                if (6'h5 == _T_168) begin
                                                                  mem_5 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h5 == _T_163) begin
                                                                    mem_5 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h5 == _T_158) begin
                                                                      mem_5 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h5 == _T_153) begin
                                                                        mem_5 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h6 == wPos) begin
            mem_6 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h6 == _T_308) begin
                mem_6 <= _GEN_31;
              end else begin
                if (6'h6 == _T_303) begin
                  mem_6 <= _GEN_30;
                end else begin
                  if (6'h6 == _T_298) begin
                    mem_6 <= _GEN_29;
                  end else begin
                    if (6'h6 == _T_293) begin
                      mem_6 <= _GEN_28;
                    end else begin
                      if (6'h6 == _T_288) begin
                        mem_6 <= _GEN_27;
                      end else begin
                        if (6'h6 == _T_283) begin
                          mem_6 <= _GEN_26;
                        end else begin
                          if (6'h6 == _T_278) begin
                            mem_6 <= _GEN_25;
                          end else begin
                            if (6'h6 == _T_273) begin
                              mem_6 <= _GEN_24;
                            end else begin
                              if (6'h6 == _T_268) begin
                                mem_6 <= _GEN_23;
                              end else begin
                                if (6'h6 == _T_263) begin
                                  mem_6 <= _GEN_22;
                                end else begin
                                  if (6'h6 == _T_258) begin
                                    mem_6 <= _GEN_21;
                                  end else begin
                                    if (6'h6 == _T_253) begin
                                      mem_6 <= _GEN_20;
                                    end else begin
                                      if (6'h6 == _T_248) begin
                                        mem_6 <= _GEN_19;
                                      end else begin
                                        if (6'h6 == _T_243) begin
                                          mem_6 <= _GEN_18;
                                        end else begin
                                          if (6'h6 == _T_238) begin
                                            mem_6 <= _GEN_17;
                                          end else begin
                                            if (6'h6 == _T_233) begin
                                              mem_6 <= _GEN_16;
                                            end else begin
                                              if (6'h6 == _T_228) begin
                                                mem_6 <= _GEN_15;
                                              end else begin
                                                if (6'h6 == _T_223) begin
                                                  mem_6 <= _GEN_14;
                                                end else begin
                                                  if (6'h6 == _T_218) begin
                                                    mem_6 <= _GEN_13;
                                                  end else begin
                                                    if (6'h6 == _T_213) begin
                                                      mem_6 <= _GEN_12;
                                                    end else begin
                                                      if (6'h6 == _T_208) begin
                                                        mem_6 <= _GEN_11;
                                                      end else begin
                                                        if (6'h6 == _T_203) begin
                                                          mem_6 <= _GEN_10;
                                                        end else begin
                                                          if (6'h6 == _T_198) begin
                                                            mem_6 <= _GEN_9;
                                                          end else begin
                                                            if (6'h6 == _T_193) begin
                                                              mem_6 <= _GEN_8;
                                                            end else begin
                                                              if (6'h6 == _T_188) begin
                                                                mem_6 <= _GEN_7;
                                                              end else begin
                                                                if (6'h6 == _T_183) begin
                                                                  mem_6 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h6 == _T_178) begin
                                                                    mem_6 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h6 == _T_173) begin
                                                                      mem_6 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h6 == _T_168) begin
                                                                        mem_6 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h6 == _T_163) begin
                                                                          mem_6 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h6 == _T_158) begin
                                                                            mem_6 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h6 == _T_153) begin
                                                                              mem_6 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h6 == _T_308) begin
              mem_6 <= _GEN_31;
            end else begin
              if (6'h6 == _T_303) begin
                mem_6 <= _GEN_30;
              end else begin
                if (6'h6 == _T_298) begin
                  mem_6 <= _GEN_29;
                end else begin
                  if (6'h6 == _T_293) begin
                    mem_6 <= _GEN_28;
                  end else begin
                    if (6'h6 == _T_288) begin
                      mem_6 <= _GEN_27;
                    end else begin
                      if (6'h6 == _T_283) begin
                        mem_6 <= _GEN_26;
                      end else begin
                        if (6'h6 == _T_278) begin
                          mem_6 <= _GEN_25;
                        end else begin
                          if (6'h6 == _T_273) begin
                            mem_6 <= _GEN_24;
                          end else begin
                            if (6'h6 == _T_268) begin
                              mem_6 <= _GEN_23;
                            end else begin
                              if (6'h6 == _T_263) begin
                                mem_6 <= _GEN_22;
                              end else begin
                                if (6'h6 == _T_258) begin
                                  mem_6 <= _GEN_21;
                                end else begin
                                  if (6'h6 == _T_253) begin
                                    mem_6 <= _GEN_20;
                                  end else begin
                                    if (6'h6 == _T_248) begin
                                      mem_6 <= _GEN_19;
                                    end else begin
                                      if (6'h6 == _T_243) begin
                                        mem_6 <= _GEN_18;
                                      end else begin
                                        if (6'h6 == _T_238) begin
                                          mem_6 <= _GEN_17;
                                        end else begin
                                          if (6'h6 == _T_233) begin
                                            mem_6 <= _GEN_16;
                                          end else begin
                                            if (6'h6 == _T_228) begin
                                              mem_6 <= _GEN_15;
                                            end else begin
                                              if (6'h6 == _T_223) begin
                                                mem_6 <= _GEN_14;
                                              end else begin
                                                if (6'h6 == _T_218) begin
                                                  mem_6 <= _GEN_13;
                                                end else begin
                                                  if (6'h6 == _T_213) begin
                                                    mem_6 <= _GEN_12;
                                                  end else begin
                                                    if (6'h6 == _T_208) begin
                                                      mem_6 <= _GEN_11;
                                                    end else begin
                                                      if (6'h6 == _T_203) begin
                                                        mem_6 <= _GEN_10;
                                                      end else begin
                                                        if (6'h6 == _T_198) begin
                                                          mem_6 <= _GEN_9;
                                                        end else begin
                                                          if (6'h6 == _T_193) begin
                                                            mem_6 <= _GEN_8;
                                                          end else begin
                                                            if (6'h6 == _T_188) begin
                                                              mem_6 <= _GEN_7;
                                                            end else begin
                                                              if (6'h6 == _T_183) begin
                                                                mem_6 <= _GEN_6;
                                                              end else begin
                                                                if (6'h6 == _T_178) begin
                                                                  mem_6 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h6 == _T_173) begin
                                                                    mem_6 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h6 == _T_168) begin
                                                                      mem_6 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h6 == _T_163) begin
                                                                        mem_6 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h6 == _T_158) begin
                                                                          mem_6 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h6 == _T_153) begin
                                                                            mem_6 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h6 == _T_308) begin
            mem_6 <= _GEN_31;
          end else begin
            if (6'h6 == _T_303) begin
              mem_6 <= _GEN_30;
            end else begin
              if (6'h6 == _T_298) begin
                mem_6 <= _GEN_29;
              end else begin
                if (6'h6 == _T_293) begin
                  mem_6 <= _GEN_28;
                end else begin
                  if (6'h6 == _T_288) begin
                    mem_6 <= _GEN_27;
                  end else begin
                    if (6'h6 == _T_283) begin
                      mem_6 <= _GEN_26;
                    end else begin
                      if (6'h6 == _T_278) begin
                        mem_6 <= _GEN_25;
                      end else begin
                        if (6'h6 == _T_273) begin
                          mem_6 <= _GEN_24;
                        end else begin
                          if (6'h6 == _T_268) begin
                            mem_6 <= _GEN_23;
                          end else begin
                            if (6'h6 == _T_263) begin
                              mem_6 <= _GEN_22;
                            end else begin
                              if (6'h6 == _T_258) begin
                                mem_6 <= _GEN_21;
                              end else begin
                                if (6'h6 == _T_253) begin
                                  mem_6 <= _GEN_20;
                                end else begin
                                  if (6'h6 == _T_248) begin
                                    mem_6 <= _GEN_19;
                                  end else begin
                                    if (6'h6 == _T_243) begin
                                      mem_6 <= _GEN_18;
                                    end else begin
                                      if (6'h6 == _T_238) begin
                                        mem_6 <= _GEN_17;
                                      end else begin
                                        if (6'h6 == _T_233) begin
                                          mem_6 <= _GEN_16;
                                        end else begin
                                          if (6'h6 == _T_228) begin
                                            mem_6 <= _GEN_15;
                                          end else begin
                                            if (6'h6 == _T_223) begin
                                              mem_6 <= _GEN_14;
                                            end else begin
                                              if (6'h6 == _T_218) begin
                                                mem_6 <= _GEN_13;
                                              end else begin
                                                if (6'h6 == _T_213) begin
                                                  mem_6 <= _GEN_12;
                                                end else begin
                                                  if (6'h6 == _T_208) begin
                                                    mem_6 <= _GEN_11;
                                                  end else begin
                                                    if (6'h6 == _T_203) begin
                                                      mem_6 <= _GEN_10;
                                                    end else begin
                                                      if (6'h6 == _T_198) begin
                                                        mem_6 <= _GEN_9;
                                                      end else begin
                                                        if (6'h6 == _T_193) begin
                                                          mem_6 <= _GEN_8;
                                                        end else begin
                                                          if (6'h6 == _T_188) begin
                                                            mem_6 <= _GEN_7;
                                                          end else begin
                                                            if (6'h6 == _T_183) begin
                                                              mem_6 <= _GEN_6;
                                                            end else begin
                                                              if (6'h6 == _T_178) begin
                                                                mem_6 <= _GEN_5;
                                                              end else begin
                                                                if (6'h6 == _T_173) begin
                                                                  mem_6 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h6 == _T_168) begin
                                                                    mem_6 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h6 == _T_163) begin
                                                                      mem_6 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h6 == _T_158) begin
                                                                        mem_6 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h6 == _T_153) begin
                                                                          mem_6 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h6 == _T_308) begin
          mem_6 <= _GEN_31;
        end else begin
          if (6'h6 == _T_303) begin
            mem_6 <= _GEN_30;
          end else begin
            if (6'h6 == _T_298) begin
              mem_6 <= _GEN_29;
            end else begin
              if (6'h6 == _T_293) begin
                mem_6 <= _GEN_28;
              end else begin
                if (6'h6 == _T_288) begin
                  mem_6 <= _GEN_27;
                end else begin
                  if (6'h6 == _T_283) begin
                    mem_6 <= _GEN_26;
                  end else begin
                    if (6'h6 == _T_278) begin
                      mem_6 <= _GEN_25;
                    end else begin
                      if (6'h6 == _T_273) begin
                        mem_6 <= _GEN_24;
                      end else begin
                        if (6'h6 == _T_268) begin
                          mem_6 <= _GEN_23;
                        end else begin
                          if (6'h6 == _T_263) begin
                            mem_6 <= _GEN_22;
                          end else begin
                            if (6'h6 == _T_258) begin
                              mem_6 <= _GEN_21;
                            end else begin
                              if (6'h6 == _T_253) begin
                                mem_6 <= _GEN_20;
                              end else begin
                                if (6'h6 == _T_248) begin
                                  mem_6 <= _GEN_19;
                                end else begin
                                  if (6'h6 == _T_243) begin
                                    mem_6 <= _GEN_18;
                                  end else begin
                                    if (6'h6 == _T_238) begin
                                      mem_6 <= _GEN_17;
                                    end else begin
                                      if (6'h6 == _T_233) begin
                                        mem_6 <= _GEN_16;
                                      end else begin
                                        if (6'h6 == _T_228) begin
                                          mem_6 <= _GEN_15;
                                        end else begin
                                          if (6'h6 == _T_223) begin
                                            mem_6 <= _GEN_14;
                                          end else begin
                                            if (6'h6 == _T_218) begin
                                              mem_6 <= _GEN_13;
                                            end else begin
                                              if (6'h6 == _T_213) begin
                                                mem_6 <= _GEN_12;
                                              end else begin
                                                if (6'h6 == _T_208) begin
                                                  mem_6 <= _GEN_11;
                                                end else begin
                                                  if (6'h6 == _T_203) begin
                                                    mem_6 <= _GEN_10;
                                                  end else begin
                                                    if (6'h6 == _T_198) begin
                                                      mem_6 <= _GEN_9;
                                                    end else begin
                                                      if (6'h6 == _T_193) begin
                                                        mem_6 <= _GEN_8;
                                                      end else begin
                                                        if (6'h6 == _T_188) begin
                                                          mem_6 <= _GEN_7;
                                                        end else begin
                                                          if (6'h6 == _T_183) begin
                                                            mem_6 <= _GEN_6;
                                                          end else begin
                                                            if (6'h6 == _T_178) begin
                                                              mem_6 <= _GEN_5;
                                                            end else begin
                                                              if (6'h6 == _T_173) begin
                                                                mem_6 <= _GEN_4;
                                                              end else begin
                                                                if (6'h6 == _T_168) begin
                                                                  mem_6 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h6 == _T_163) begin
                                                                    mem_6 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h6 == _T_158) begin
                                                                      mem_6 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h6 == _T_153) begin
                                                                        mem_6 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h7 == wPos) begin
            mem_7 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h7 == _T_308) begin
                mem_7 <= _GEN_31;
              end else begin
                if (6'h7 == _T_303) begin
                  mem_7 <= _GEN_30;
                end else begin
                  if (6'h7 == _T_298) begin
                    mem_7 <= _GEN_29;
                  end else begin
                    if (6'h7 == _T_293) begin
                      mem_7 <= _GEN_28;
                    end else begin
                      if (6'h7 == _T_288) begin
                        mem_7 <= _GEN_27;
                      end else begin
                        if (6'h7 == _T_283) begin
                          mem_7 <= _GEN_26;
                        end else begin
                          if (6'h7 == _T_278) begin
                            mem_7 <= _GEN_25;
                          end else begin
                            if (6'h7 == _T_273) begin
                              mem_7 <= _GEN_24;
                            end else begin
                              if (6'h7 == _T_268) begin
                                mem_7 <= _GEN_23;
                              end else begin
                                if (6'h7 == _T_263) begin
                                  mem_7 <= _GEN_22;
                                end else begin
                                  if (6'h7 == _T_258) begin
                                    mem_7 <= _GEN_21;
                                  end else begin
                                    if (6'h7 == _T_253) begin
                                      mem_7 <= _GEN_20;
                                    end else begin
                                      if (6'h7 == _T_248) begin
                                        mem_7 <= _GEN_19;
                                      end else begin
                                        if (6'h7 == _T_243) begin
                                          mem_7 <= _GEN_18;
                                        end else begin
                                          if (6'h7 == _T_238) begin
                                            mem_7 <= _GEN_17;
                                          end else begin
                                            if (6'h7 == _T_233) begin
                                              mem_7 <= _GEN_16;
                                            end else begin
                                              if (6'h7 == _T_228) begin
                                                mem_7 <= _GEN_15;
                                              end else begin
                                                if (6'h7 == _T_223) begin
                                                  mem_7 <= _GEN_14;
                                                end else begin
                                                  if (6'h7 == _T_218) begin
                                                    mem_7 <= _GEN_13;
                                                  end else begin
                                                    if (6'h7 == _T_213) begin
                                                      mem_7 <= _GEN_12;
                                                    end else begin
                                                      if (6'h7 == _T_208) begin
                                                        mem_7 <= _GEN_11;
                                                      end else begin
                                                        if (6'h7 == _T_203) begin
                                                          mem_7 <= _GEN_10;
                                                        end else begin
                                                          if (6'h7 == _T_198) begin
                                                            mem_7 <= _GEN_9;
                                                          end else begin
                                                            if (6'h7 == _T_193) begin
                                                              mem_7 <= _GEN_8;
                                                            end else begin
                                                              if (6'h7 == _T_188) begin
                                                                mem_7 <= _GEN_7;
                                                              end else begin
                                                                if (6'h7 == _T_183) begin
                                                                  mem_7 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h7 == _T_178) begin
                                                                    mem_7 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h7 == _T_173) begin
                                                                      mem_7 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h7 == _T_168) begin
                                                                        mem_7 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h7 == _T_163) begin
                                                                          mem_7 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h7 == _T_158) begin
                                                                            mem_7 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h7 == _T_153) begin
                                                                              mem_7 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h7 == _T_308) begin
              mem_7 <= _GEN_31;
            end else begin
              if (6'h7 == _T_303) begin
                mem_7 <= _GEN_30;
              end else begin
                if (6'h7 == _T_298) begin
                  mem_7 <= _GEN_29;
                end else begin
                  if (6'h7 == _T_293) begin
                    mem_7 <= _GEN_28;
                  end else begin
                    if (6'h7 == _T_288) begin
                      mem_7 <= _GEN_27;
                    end else begin
                      if (6'h7 == _T_283) begin
                        mem_7 <= _GEN_26;
                      end else begin
                        if (6'h7 == _T_278) begin
                          mem_7 <= _GEN_25;
                        end else begin
                          if (6'h7 == _T_273) begin
                            mem_7 <= _GEN_24;
                          end else begin
                            if (6'h7 == _T_268) begin
                              mem_7 <= _GEN_23;
                            end else begin
                              if (6'h7 == _T_263) begin
                                mem_7 <= _GEN_22;
                              end else begin
                                if (6'h7 == _T_258) begin
                                  mem_7 <= _GEN_21;
                                end else begin
                                  if (6'h7 == _T_253) begin
                                    mem_7 <= _GEN_20;
                                  end else begin
                                    if (6'h7 == _T_248) begin
                                      mem_7 <= _GEN_19;
                                    end else begin
                                      if (6'h7 == _T_243) begin
                                        mem_7 <= _GEN_18;
                                      end else begin
                                        if (6'h7 == _T_238) begin
                                          mem_7 <= _GEN_17;
                                        end else begin
                                          if (6'h7 == _T_233) begin
                                            mem_7 <= _GEN_16;
                                          end else begin
                                            if (6'h7 == _T_228) begin
                                              mem_7 <= _GEN_15;
                                            end else begin
                                              if (6'h7 == _T_223) begin
                                                mem_7 <= _GEN_14;
                                              end else begin
                                                if (6'h7 == _T_218) begin
                                                  mem_7 <= _GEN_13;
                                                end else begin
                                                  if (6'h7 == _T_213) begin
                                                    mem_7 <= _GEN_12;
                                                  end else begin
                                                    if (6'h7 == _T_208) begin
                                                      mem_7 <= _GEN_11;
                                                    end else begin
                                                      if (6'h7 == _T_203) begin
                                                        mem_7 <= _GEN_10;
                                                      end else begin
                                                        if (6'h7 == _T_198) begin
                                                          mem_7 <= _GEN_9;
                                                        end else begin
                                                          if (6'h7 == _T_193) begin
                                                            mem_7 <= _GEN_8;
                                                          end else begin
                                                            if (6'h7 == _T_188) begin
                                                              mem_7 <= _GEN_7;
                                                            end else begin
                                                              if (6'h7 == _T_183) begin
                                                                mem_7 <= _GEN_6;
                                                              end else begin
                                                                if (6'h7 == _T_178) begin
                                                                  mem_7 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h7 == _T_173) begin
                                                                    mem_7 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h7 == _T_168) begin
                                                                      mem_7 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h7 == _T_163) begin
                                                                        mem_7 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h7 == _T_158) begin
                                                                          mem_7 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h7 == _T_153) begin
                                                                            mem_7 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h7 == _T_308) begin
            mem_7 <= _GEN_31;
          end else begin
            if (6'h7 == _T_303) begin
              mem_7 <= _GEN_30;
            end else begin
              if (6'h7 == _T_298) begin
                mem_7 <= _GEN_29;
              end else begin
                if (6'h7 == _T_293) begin
                  mem_7 <= _GEN_28;
                end else begin
                  if (6'h7 == _T_288) begin
                    mem_7 <= _GEN_27;
                  end else begin
                    if (6'h7 == _T_283) begin
                      mem_7 <= _GEN_26;
                    end else begin
                      if (6'h7 == _T_278) begin
                        mem_7 <= _GEN_25;
                      end else begin
                        if (6'h7 == _T_273) begin
                          mem_7 <= _GEN_24;
                        end else begin
                          if (6'h7 == _T_268) begin
                            mem_7 <= _GEN_23;
                          end else begin
                            if (6'h7 == _T_263) begin
                              mem_7 <= _GEN_22;
                            end else begin
                              if (6'h7 == _T_258) begin
                                mem_7 <= _GEN_21;
                              end else begin
                                if (6'h7 == _T_253) begin
                                  mem_7 <= _GEN_20;
                                end else begin
                                  if (6'h7 == _T_248) begin
                                    mem_7 <= _GEN_19;
                                  end else begin
                                    if (6'h7 == _T_243) begin
                                      mem_7 <= _GEN_18;
                                    end else begin
                                      if (6'h7 == _T_238) begin
                                        mem_7 <= _GEN_17;
                                      end else begin
                                        if (6'h7 == _T_233) begin
                                          mem_7 <= _GEN_16;
                                        end else begin
                                          if (6'h7 == _T_228) begin
                                            mem_7 <= _GEN_15;
                                          end else begin
                                            if (6'h7 == _T_223) begin
                                              mem_7 <= _GEN_14;
                                            end else begin
                                              if (6'h7 == _T_218) begin
                                                mem_7 <= _GEN_13;
                                              end else begin
                                                if (6'h7 == _T_213) begin
                                                  mem_7 <= _GEN_12;
                                                end else begin
                                                  if (6'h7 == _T_208) begin
                                                    mem_7 <= _GEN_11;
                                                  end else begin
                                                    if (6'h7 == _T_203) begin
                                                      mem_7 <= _GEN_10;
                                                    end else begin
                                                      if (6'h7 == _T_198) begin
                                                        mem_7 <= _GEN_9;
                                                      end else begin
                                                        if (6'h7 == _T_193) begin
                                                          mem_7 <= _GEN_8;
                                                        end else begin
                                                          if (6'h7 == _T_188) begin
                                                            mem_7 <= _GEN_7;
                                                          end else begin
                                                            if (6'h7 == _T_183) begin
                                                              mem_7 <= _GEN_6;
                                                            end else begin
                                                              if (6'h7 == _T_178) begin
                                                                mem_7 <= _GEN_5;
                                                              end else begin
                                                                if (6'h7 == _T_173) begin
                                                                  mem_7 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h7 == _T_168) begin
                                                                    mem_7 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h7 == _T_163) begin
                                                                      mem_7 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h7 == _T_158) begin
                                                                        mem_7 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h7 == _T_153) begin
                                                                          mem_7 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h7 == _T_308) begin
          mem_7 <= _GEN_31;
        end else begin
          if (6'h7 == _T_303) begin
            mem_7 <= _GEN_30;
          end else begin
            if (6'h7 == _T_298) begin
              mem_7 <= _GEN_29;
            end else begin
              if (6'h7 == _T_293) begin
                mem_7 <= _GEN_28;
              end else begin
                if (6'h7 == _T_288) begin
                  mem_7 <= _GEN_27;
                end else begin
                  if (6'h7 == _T_283) begin
                    mem_7 <= _GEN_26;
                  end else begin
                    if (6'h7 == _T_278) begin
                      mem_7 <= _GEN_25;
                    end else begin
                      if (6'h7 == _T_273) begin
                        mem_7 <= _GEN_24;
                      end else begin
                        if (6'h7 == _T_268) begin
                          mem_7 <= _GEN_23;
                        end else begin
                          if (6'h7 == _T_263) begin
                            mem_7 <= _GEN_22;
                          end else begin
                            if (6'h7 == _T_258) begin
                              mem_7 <= _GEN_21;
                            end else begin
                              if (6'h7 == _T_253) begin
                                mem_7 <= _GEN_20;
                              end else begin
                                if (6'h7 == _T_248) begin
                                  mem_7 <= _GEN_19;
                                end else begin
                                  if (6'h7 == _T_243) begin
                                    mem_7 <= _GEN_18;
                                  end else begin
                                    if (6'h7 == _T_238) begin
                                      mem_7 <= _GEN_17;
                                    end else begin
                                      if (6'h7 == _T_233) begin
                                        mem_7 <= _GEN_16;
                                      end else begin
                                        if (6'h7 == _T_228) begin
                                          mem_7 <= _GEN_15;
                                        end else begin
                                          if (6'h7 == _T_223) begin
                                            mem_7 <= _GEN_14;
                                          end else begin
                                            if (6'h7 == _T_218) begin
                                              mem_7 <= _GEN_13;
                                            end else begin
                                              if (6'h7 == _T_213) begin
                                                mem_7 <= _GEN_12;
                                              end else begin
                                                if (6'h7 == _T_208) begin
                                                  mem_7 <= _GEN_11;
                                                end else begin
                                                  if (6'h7 == _T_203) begin
                                                    mem_7 <= _GEN_10;
                                                  end else begin
                                                    if (6'h7 == _T_198) begin
                                                      mem_7 <= _GEN_9;
                                                    end else begin
                                                      if (6'h7 == _T_193) begin
                                                        mem_7 <= _GEN_8;
                                                      end else begin
                                                        if (6'h7 == _T_188) begin
                                                          mem_7 <= _GEN_7;
                                                        end else begin
                                                          if (6'h7 == _T_183) begin
                                                            mem_7 <= _GEN_6;
                                                          end else begin
                                                            if (6'h7 == _T_178) begin
                                                              mem_7 <= _GEN_5;
                                                            end else begin
                                                              if (6'h7 == _T_173) begin
                                                                mem_7 <= _GEN_4;
                                                              end else begin
                                                                if (6'h7 == _T_168) begin
                                                                  mem_7 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h7 == _T_163) begin
                                                                    mem_7 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h7 == _T_158) begin
                                                                      mem_7 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h7 == _T_153) begin
                                                                        mem_7 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h8 == wPos) begin
            mem_8 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h8 == _T_308) begin
                mem_8 <= _GEN_31;
              end else begin
                if (6'h8 == _T_303) begin
                  mem_8 <= _GEN_30;
                end else begin
                  if (6'h8 == _T_298) begin
                    mem_8 <= _GEN_29;
                  end else begin
                    if (6'h8 == _T_293) begin
                      mem_8 <= _GEN_28;
                    end else begin
                      if (6'h8 == _T_288) begin
                        mem_8 <= _GEN_27;
                      end else begin
                        if (6'h8 == _T_283) begin
                          mem_8 <= _GEN_26;
                        end else begin
                          if (6'h8 == _T_278) begin
                            mem_8 <= _GEN_25;
                          end else begin
                            if (6'h8 == _T_273) begin
                              mem_8 <= _GEN_24;
                            end else begin
                              if (6'h8 == _T_268) begin
                                mem_8 <= _GEN_23;
                              end else begin
                                if (6'h8 == _T_263) begin
                                  mem_8 <= _GEN_22;
                                end else begin
                                  if (6'h8 == _T_258) begin
                                    mem_8 <= _GEN_21;
                                  end else begin
                                    if (6'h8 == _T_253) begin
                                      mem_8 <= _GEN_20;
                                    end else begin
                                      if (6'h8 == _T_248) begin
                                        mem_8 <= _GEN_19;
                                      end else begin
                                        if (6'h8 == _T_243) begin
                                          mem_8 <= _GEN_18;
                                        end else begin
                                          if (6'h8 == _T_238) begin
                                            mem_8 <= _GEN_17;
                                          end else begin
                                            if (6'h8 == _T_233) begin
                                              mem_8 <= _GEN_16;
                                            end else begin
                                              if (6'h8 == _T_228) begin
                                                mem_8 <= _GEN_15;
                                              end else begin
                                                if (6'h8 == _T_223) begin
                                                  mem_8 <= _GEN_14;
                                                end else begin
                                                  if (6'h8 == _T_218) begin
                                                    mem_8 <= _GEN_13;
                                                  end else begin
                                                    if (6'h8 == _T_213) begin
                                                      mem_8 <= _GEN_12;
                                                    end else begin
                                                      if (6'h8 == _T_208) begin
                                                        mem_8 <= _GEN_11;
                                                      end else begin
                                                        if (6'h8 == _T_203) begin
                                                          mem_8 <= _GEN_10;
                                                        end else begin
                                                          if (6'h8 == _T_198) begin
                                                            mem_8 <= _GEN_9;
                                                          end else begin
                                                            if (6'h8 == _T_193) begin
                                                              mem_8 <= _GEN_8;
                                                            end else begin
                                                              if (6'h8 == _T_188) begin
                                                                mem_8 <= _GEN_7;
                                                              end else begin
                                                                if (6'h8 == _T_183) begin
                                                                  mem_8 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h8 == _T_178) begin
                                                                    mem_8 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h8 == _T_173) begin
                                                                      mem_8 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h8 == _T_168) begin
                                                                        mem_8 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h8 == _T_163) begin
                                                                          mem_8 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h8 == _T_158) begin
                                                                            mem_8 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h8 == _T_153) begin
                                                                              mem_8 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h8 == _T_308) begin
              mem_8 <= _GEN_31;
            end else begin
              if (6'h8 == _T_303) begin
                mem_8 <= _GEN_30;
              end else begin
                if (6'h8 == _T_298) begin
                  mem_8 <= _GEN_29;
                end else begin
                  if (6'h8 == _T_293) begin
                    mem_8 <= _GEN_28;
                  end else begin
                    if (6'h8 == _T_288) begin
                      mem_8 <= _GEN_27;
                    end else begin
                      if (6'h8 == _T_283) begin
                        mem_8 <= _GEN_26;
                      end else begin
                        if (6'h8 == _T_278) begin
                          mem_8 <= _GEN_25;
                        end else begin
                          if (6'h8 == _T_273) begin
                            mem_8 <= _GEN_24;
                          end else begin
                            if (6'h8 == _T_268) begin
                              mem_8 <= _GEN_23;
                            end else begin
                              if (6'h8 == _T_263) begin
                                mem_8 <= _GEN_22;
                              end else begin
                                if (6'h8 == _T_258) begin
                                  mem_8 <= _GEN_21;
                                end else begin
                                  if (6'h8 == _T_253) begin
                                    mem_8 <= _GEN_20;
                                  end else begin
                                    if (6'h8 == _T_248) begin
                                      mem_8 <= _GEN_19;
                                    end else begin
                                      if (6'h8 == _T_243) begin
                                        mem_8 <= _GEN_18;
                                      end else begin
                                        if (6'h8 == _T_238) begin
                                          mem_8 <= _GEN_17;
                                        end else begin
                                          if (6'h8 == _T_233) begin
                                            mem_8 <= _GEN_16;
                                          end else begin
                                            if (6'h8 == _T_228) begin
                                              mem_8 <= _GEN_15;
                                            end else begin
                                              if (6'h8 == _T_223) begin
                                                mem_8 <= _GEN_14;
                                              end else begin
                                                if (6'h8 == _T_218) begin
                                                  mem_8 <= _GEN_13;
                                                end else begin
                                                  if (6'h8 == _T_213) begin
                                                    mem_8 <= _GEN_12;
                                                  end else begin
                                                    if (6'h8 == _T_208) begin
                                                      mem_8 <= _GEN_11;
                                                    end else begin
                                                      if (6'h8 == _T_203) begin
                                                        mem_8 <= _GEN_10;
                                                      end else begin
                                                        if (6'h8 == _T_198) begin
                                                          mem_8 <= _GEN_9;
                                                        end else begin
                                                          if (6'h8 == _T_193) begin
                                                            mem_8 <= _GEN_8;
                                                          end else begin
                                                            if (6'h8 == _T_188) begin
                                                              mem_8 <= _GEN_7;
                                                            end else begin
                                                              if (6'h8 == _T_183) begin
                                                                mem_8 <= _GEN_6;
                                                              end else begin
                                                                if (6'h8 == _T_178) begin
                                                                  mem_8 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h8 == _T_173) begin
                                                                    mem_8 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h8 == _T_168) begin
                                                                      mem_8 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h8 == _T_163) begin
                                                                        mem_8 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h8 == _T_158) begin
                                                                          mem_8 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h8 == _T_153) begin
                                                                            mem_8 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h8 == _T_308) begin
            mem_8 <= _GEN_31;
          end else begin
            if (6'h8 == _T_303) begin
              mem_8 <= _GEN_30;
            end else begin
              if (6'h8 == _T_298) begin
                mem_8 <= _GEN_29;
              end else begin
                if (6'h8 == _T_293) begin
                  mem_8 <= _GEN_28;
                end else begin
                  if (6'h8 == _T_288) begin
                    mem_8 <= _GEN_27;
                  end else begin
                    if (6'h8 == _T_283) begin
                      mem_8 <= _GEN_26;
                    end else begin
                      if (6'h8 == _T_278) begin
                        mem_8 <= _GEN_25;
                      end else begin
                        if (6'h8 == _T_273) begin
                          mem_8 <= _GEN_24;
                        end else begin
                          if (6'h8 == _T_268) begin
                            mem_8 <= _GEN_23;
                          end else begin
                            if (6'h8 == _T_263) begin
                              mem_8 <= _GEN_22;
                            end else begin
                              if (6'h8 == _T_258) begin
                                mem_8 <= _GEN_21;
                              end else begin
                                if (6'h8 == _T_253) begin
                                  mem_8 <= _GEN_20;
                                end else begin
                                  if (6'h8 == _T_248) begin
                                    mem_8 <= _GEN_19;
                                  end else begin
                                    if (6'h8 == _T_243) begin
                                      mem_8 <= _GEN_18;
                                    end else begin
                                      if (6'h8 == _T_238) begin
                                        mem_8 <= _GEN_17;
                                      end else begin
                                        if (6'h8 == _T_233) begin
                                          mem_8 <= _GEN_16;
                                        end else begin
                                          if (6'h8 == _T_228) begin
                                            mem_8 <= _GEN_15;
                                          end else begin
                                            if (6'h8 == _T_223) begin
                                              mem_8 <= _GEN_14;
                                            end else begin
                                              if (6'h8 == _T_218) begin
                                                mem_8 <= _GEN_13;
                                              end else begin
                                                if (6'h8 == _T_213) begin
                                                  mem_8 <= _GEN_12;
                                                end else begin
                                                  if (6'h8 == _T_208) begin
                                                    mem_8 <= _GEN_11;
                                                  end else begin
                                                    if (6'h8 == _T_203) begin
                                                      mem_8 <= _GEN_10;
                                                    end else begin
                                                      if (6'h8 == _T_198) begin
                                                        mem_8 <= _GEN_9;
                                                      end else begin
                                                        if (6'h8 == _T_193) begin
                                                          mem_8 <= _GEN_8;
                                                        end else begin
                                                          if (6'h8 == _T_188) begin
                                                            mem_8 <= _GEN_7;
                                                          end else begin
                                                            if (6'h8 == _T_183) begin
                                                              mem_8 <= _GEN_6;
                                                            end else begin
                                                              if (6'h8 == _T_178) begin
                                                                mem_8 <= _GEN_5;
                                                              end else begin
                                                                if (6'h8 == _T_173) begin
                                                                  mem_8 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h8 == _T_168) begin
                                                                    mem_8 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h8 == _T_163) begin
                                                                      mem_8 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h8 == _T_158) begin
                                                                        mem_8 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h8 == _T_153) begin
                                                                          mem_8 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h8 == _T_308) begin
          mem_8 <= _GEN_31;
        end else begin
          if (6'h8 == _T_303) begin
            mem_8 <= _GEN_30;
          end else begin
            if (6'h8 == _T_298) begin
              mem_8 <= _GEN_29;
            end else begin
              if (6'h8 == _T_293) begin
                mem_8 <= _GEN_28;
              end else begin
                if (6'h8 == _T_288) begin
                  mem_8 <= _GEN_27;
                end else begin
                  if (6'h8 == _T_283) begin
                    mem_8 <= _GEN_26;
                  end else begin
                    if (6'h8 == _T_278) begin
                      mem_8 <= _GEN_25;
                    end else begin
                      if (6'h8 == _T_273) begin
                        mem_8 <= _GEN_24;
                      end else begin
                        if (6'h8 == _T_268) begin
                          mem_8 <= _GEN_23;
                        end else begin
                          if (6'h8 == _T_263) begin
                            mem_8 <= _GEN_22;
                          end else begin
                            if (6'h8 == _T_258) begin
                              mem_8 <= _GEN_21;
                            end else begin
                              if (6'h8 == _T_253) begin
                                mem_8 <= _GEN_20;
                              end else begin
                                if (6'h8 == _T_248) begin
                                  mem_8 <= _GEN_19;
                                end else begin
                                  if (6'h8 == _T_243) begin
                                    mem_8 <= _GEN_18;
                                  end else begin
                                    if (6'h8 == _T_238) begin
                                      mem_8 <= _GEN_17;
                                    end else begin
                                      if (6'h8 == _T_233) begin
                                        mem_8 <= _GEN_16;
                                      end else begin
                                        if (6'h8 == _T_228) begin
                                          mem_8 <= _GEN_15;
                                        end else begin
                                          if (6'h8 == _T_223) begin
                                            mem_8 <= _GEN_14;
                                          end else begin
                                            if (6'h8 == _T_218) begin
                                              mem_8 <= _GEN_13;
                                            end else begin
                                              if (6'h8 == _T_213) begin
                                                mem_8 <= _GEN_12;
                                              end else begin
                                                if (6'h8 == _T_208) begin
                                                  mem_8 <= _GEN_11;
                                                end else begin
                                                  if (6'h8 == _T_203) begin
                                                    mem_8 <= _GEN_10;
                                                  end else begin
                                                    if (6'h8 == _T_198) begin
                                                      mem_8 <= _GEN_9;
                                                    end else begin
                                                      if (6'h8 == _T_193) begin
                                                        mem_8 <= _GEN_8;
                                                      end else begin
                                                        if (6'h8 == _T_188) begin
                                                          mem_8 <= _GEN_7;
                                                        end else begin
                                                          if (6'h8 == _T_183) begin
                                                            mem_8 <= _GEN_6;
                                                          end else begin
                                                            if (6'h8 == _T_178) begin
                                                              mem_8 <= _GEN_5;
                                                            end else begin
                                                              if (6'h8 == _T_173) begin
                                                                mem_8 <= _GEN_4;
                                                              end else begin
                                                                if (6'h8 == _T_168) begin
                                                                  mem_8 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h8 == _T_163) begin
                                                                    mem_8 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h8 == _T_158) begin
                                                                      mem_8 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h8 == _T_153) begin
                                                                        mem_8 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h9 == wPos) begin
            mem_9 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h9 == _T_308) begin
                mem_9 <= _GEN_31;
              end else begin
                if (6'h9 == _T_303) begin
                  mem_9 <= _GEN_30;
                end else begin
                  if (6'h9 == _T_298) begin
                    mem_9 <= _GEN_29;
                  end else begin
                    if (6'h9 == _T_293) begin
                      mem_9 <= _GEN_28;
                    end else begin
                      if (6'h9 == _T_288) begin
                        mem_9 <= _GEN_27;
                      end else begin
                        if (6'h9 == _T_283) begin
                          mem_9 <= _GEN_26;
                        end else begin
                          if (6'h9 == _T_278) begin
                            mem_9 <= _GEN_25;
                          end else begin
                            if (6'h9 == _T_273) begin
                              mem_9 <= _GEN_24;
                            end else begin
                              if (6'h9 == _T_268) begin
                                mem_9 <= _GEN_23;
                              end else begin
                                if (6'h9 == _T_263) begin
                                  mem_9 <= _GEN_22;
                                end else begin
                                  if (6'h9 == _T_258) begin
                                    mem_9 <= _GEN_21;
                                  end else begin
                                    if (6'h9 == _T_253) begin
                                      mem_9 <= _GEN_20;
                                    end else begin
                                      if (6'h9 == _T_248) begin
                                        mem_9 <= _GEN_19;
                                      end else begin
                                        if (6'h9 == _T_243) begin
                                          mem_9 <= _GEN_18;
                                        end else begin
                                          if (6'h9 == _T_238) begin
                                            mem_9 <= _GEN_17;
                                          end else begin
                                            if (6'h9 == _T_233) begin
                                              mem_9 <= _GEN_16;
                                            end else begin
                                              if (6'h9 == _T_228) begin
                                                mem_9 <= _GEN_15;
                                              end else begin
                                                if (6'h9 == _T_223) begin
                                                  mem_9 <= _GEN_14;
                                                end else begin
                                                  if (6'h9 == _T_218) begin
                                                    mem_9 <= _GEN_13;
                                                  end else begin
                                                    if (6'h9 == _T_213) begin
                                                      mem_9 <= _GEN_12;
                                                    end else begin
                                                      if (6'h9 == _T_208) begin
                                                        mem_9 <= _GEN_11;
                                                      end else begin
                                                        if (6'h9 == _T_203) begin
                                                          mem_9 <= _GEN_10;
                                                        end else begin
                                                          if (6'h9 == _T_198) begin
                                                            mem_9 <= _GEN_9;
                                                          end else begin
                                                            if (6'h9 == _T_193) begin
                                                              mem_9 <= _GEN_8;
                                                            end else begin
                                                              if (6'h9 == _T_188) begin
                                                                mem_9 <= _GEN_7;
                                                              end else begin
                                                                if (6'h9 == _T_183) begin
                                                                  mem_9 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h9 == _T_178) begin
                                                                    mem_9 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h9 == _T_173) begin
                                                                      mem_9 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h9 == _T_168) begin
                                                                        mem_9 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h9 == _T_163) begin
                                                                          mem_9 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h9 == _T_158) begin
                                                                            mem_9 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h9 == _T_153) begin
                                                                              mem_9 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h9 == _T_308) begin
              mem_9 <= _GEN_31;
            end else begin
              if (6'h9 == _T_303) begin
                mem_9 <= _GEN_30;
              end else begin
                if (6'h9 == _T_298) begin
                  mem_9 <= _GEN_29;
                end else begin
                  if (6'h9 == _T_293) begin
                    mem_9 <= _GEN_28;
                  end else begin
                    if (6'h9 == _T_288) begin
                      mem_9 <= _GEN_27;
                    end else begin
                      if (6'h9 == _T_283) begin
                        mem_9 <= _GEN_26;
                      end else begin
                        if (6'h9 == _T_278) begin
                          mem_9 <= _GEN_25;
                        end else begin
                          if (6'h9 == _T_273) begin
                            mem_9 <= _GEN_24;
                          end else begin
                            if (6'h9 == _T_268) begin
                              mem_9 <= _GEN_23;
                            end else begin
                              if (6'h9 == _T_263) begin
                                mem_9 <= _GEN_22;
                              end else begin
                                if (6'h9 == _T_258) begin
                                  mem_9 <= _GEN_21;
                                end else begin
                                  if (6'h9 == _T_253) begin
                                    mem_9 <= _GEN_20;
                                  end else begin
                                    if (6'h9 == _T_248) begin
                                      mem_9 <= _GEN_19;
                                    end else begin
                                      if (6'h9 == _T_243) begin
                                        mem_9 <= _GEN_18;
                                      end else begin
                                        if (6'h9 == _T_238) begin
                                          mem_9 <= _GEN_17;
                                        end else begin
                                          if (6'h9 == _T_233) begin
                                            mem_9 <= _GEN_16;
                                          end else begin
                                            if (6'h9 == _T_228) begin
                                              mem_9 <= _GEN_15;
                                            end else begin
                                              if (6'h9 == _T_223) begin
                                                mem_9 <= _GEN_14;
                                              end else begin
                                                if (6'h9 == _T_218) begin
                                                  mem_9 <= _GEN_13;
                                                end else begin
                                                  if (6'h9 == _T_213) begin
                                                    mem_9 <= _GEN_12;
                                                  end else begin
                                                    if (6'h9 == _T_208) begin
                                                      mem_9 <= _GEN_11;
                                                    end else begin
                                                      if (6'h9 == _T_203) begin
                                                        mem_9 <= _GEN_10;
                                                      end else begin
                                                        if (6'h9 == _T_198) begin
                                                          mem_9 <= _GEN_9;
                                                        end else begin
                                                          if (6'h9 == _T_193) begin
                                                            mem_9 <= _GEN_8;
                                                          end else begin
                                                            if (6'h9 == _T_188) begin
                                                              mem_9 <= _GEN_7;
                                                            end else begin
                                                              if (6'h9 == _T_183) begin
                                                                mem_9 <= _GEN_6;
                                                              end else begin
                                                                if (6'h9 == _T_178) begin
                                                                  mem_9 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h9 == _T_173) begin
                                                                    mem_9 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h9 == _T_168) begin
                                                                      mem_9 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h9 == _T_163) begin
                                                                        mem_9 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h9 == _T_158) begin
                                                                          mem_9 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h9 == _T_153) begin
                                                                            mem_9 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h9 == _T_308) begin
            mem_9 <= _GEN_31;
          end else begin
            if (6'h9 == _T_303) begin
              mem_9 <= _GEN_30;
            end else begin
              if (6'h9 == _T_298) begin
                mem_9 <= _GEN_29;
              end else begin
                if (6'h9 == _T_293) begin
                  mem_9 <= _GEN_28;
                end else begin
                  if (6'h9 == _T_288) begin
                    mem_9 <= _GEN_27;
                  end else begin
                    if (6'h9 == _T_283) begin
                      mem_9 <= _GEN_26;
                    end else begin
                      if (6'h9 == _T_278) begin
                        mem_9 <= _GEN_25;
                      end else begin
                        if (6'h9 == _T_273) begin
                          mem_9 <= _GEN_24;
                        end else begin
                          if (6'h9 == _T_268) begin
                            mem_9 <= _GEN_23;
                          end else begin
                            if (6'h9 == _T_263) begin
                              mem_9 <= _GEN_22;
                            end else begin
                              if (6'h9 == _T_258) begin
                                mem_9 <= _GEN_21;
                              end else begin
                                if (6'h9 == _T_253) begin
                                  mem_9 <= _GEN_20;
                                end else begin
                                  if (6'h9 == _T_248) begin
                                    mem_9 <= _GEN_19;
                                  end else begin
                                    if (6'h9 == _T_243) begin
                                      mem_9 <= _GEN_18;
                                    end else begin
                                      if (6'h9 == _T_238) begin
                                        mem_9 <= _GEN_17;
                                      end else begin
                                        if (6'h9 == _T_233) begin
                                          mem_9 <= _GEN_16;
                                        end else begin
                                          if (6'h9 == _T_228) begin
                                            mem_9 <= _GEN_15;
                                          end else begin
                                            if (6'h9 == _T_223) begin
                                              mem_9 <= _GEN_14;
                                            end else begin
                                              if (6'h9 == _T_218) begin
                                                mem_9 <= _GEN_13;
                                              end else begin
                                                if (6'h9 == _T_213) begin
                                                  mem_9 <= _GEN_12;
                                                end else begin
                                                  if (6'h9 == _T_208) begin
                                                    mem_9 <= _GEN_11;
                                                  end else begin
                                                    if (6'h9 == _T_203) begin
                                                      mem_9 <= _GEN_10;
                                                    end else begin
                                                      if (6'h9 == _T_198) begin
                                                        mem_9 <= _GEN_9;
                                                      end else begin
                                                        if (6'h9 == _T_193) begin
                                                          mem_9 <= _GEN_8;
                                                        end else begin
                                                          if (6'h9 == _T_188) begin
                                                            mem_9 <= _GEN_7;
                                                          end else begin
                                                            if (6'h9 == _T_183) begin
                                                              mem_9 <= _GEN_6;
                                                            end else begin
                                                              if (6'h9 == _T_178) begin
                                                                mem_9 <= _GEN_5;
                                                              end else begin
                                                                if (6'h9 == _T_173) begin
                                                                  mem_9 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h9 == _T_168) begin
                                                                    mem_9 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h9 == _T_163) begin
                                                                      mem_9 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h9 == _T_158) begin
                                                                        mem_9 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h9 == _T_153) begin
                                                                          mem_9 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h9 == _T_308) begin
          mem_9 <= _GEN_31;
        end else begin
          if (6'h9 == _T_303) begin
            mem_9 <= _GEN_30;
          end else begin
            if (6'h9 == _T_298) begin
              mem_9 <= _GEN_29;
            end else begin
              if (6'h9 == _T_293) begin
                mem_9 <= _GEN_28;
              end else begin
                if (6'h9 == _T_288) begin
                  mem_9 <= _GEN_27;
                end else begin
                  if (6'h9 == _T_283) begin
                    mem_9 <= _GEN_26;
                  end else begin
                    if (6'h9 == _T_278) begin
                      mem_9 <= _GEN_25;
                    end else begin
                      if (6'h9 == _T_273) begin
                        mem_9 <= _GEN_24;
                      end else begin
                        if (6'h9 == _T_268) begin
                          mem_9 <= _GEN_23;
                        end else begin
                          if (6'h9 == _T_263) begin
                            mem_9 <= _GEN_22;
                          end else begin
                            if (6'h9 == _T_258) begin
                              mem_9 <= _GEN_21;
                            end else begin
                              if (6'h9 == _T_253) begin
                                mem_9 <= _GEN_20;
                              end else begin
                                if (6'h9 == _T_248) begin
                                  mem_9 <= _GEN_19;
                                end else begin
                                  if (6'h9 == _T_243) begin
                                    mem_9 <= _GEN_18;
                                  end else begin
                                    if (6'h9 == _T_238) begin
                                      mem_9 <= _GEN_17;
                                    end else begin
                                      if (6'h9 == _T_233) begin
                                        mem_9 <= _GEN_16;
                                      end else begin
                                        if (6'h9 == _T_228) begin
                                          mem_9 <= _GEN_15;
                                        end else begin
                                          if (6'h9 == _T_223) begin
                                            mem_9 <= _GEN_14;
                                          end else begin
                                            if (6'h9 == _T_218) begin
                                              mem_9 <= _GEN_13;
                                            end else begin
                                              if (6'h9 == _T_213) begin
                                                mem_9 <= _GEN_12;
                                              end else begin
                                                if (6'h9 == _T_208) begin
                                                  mem_9 <= _GEN_11;
                                                end else begin
                                                  if (6'h9 == _T_203) begin
                                                    mem_9 <= _GEN_10;
                                                  end else begin
                                                    if (6'h9 == _T_198) begin
                                                      mem_9 <= _GEN_9;
                                                    end else begin
                                                      if (6'h9 == _T_193) begin
                                                        mem_9 <= _GEN_8;
                                                      end else begin
                                                        if (6'h9 == _T_188) begin
                                                          mem_9 <= _GEN_7;
                                                        end else begin
                                                          if (6'h9 == _T_183) begin
                                                            mem_9 <= _GEN_6;
                                                          end else begin
                                                            if (6'h9 == _T_178) begin
                                                              mem_9 <= _GEN_5;
                                                            end else begin
                                                              if (6'h9 == _T_173) begin
                                                                mem_9 <= _GEN_4;
                                                              end else begin
                                                                if (6'h9 == _T_168) begin
                                                                  mem_9 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h9 == _T_163) begin
                                                                    mem_9 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h9 == _T_158) begin
                                                                      mem_9 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h9 == _T_153) begin
                                                                        mem_9 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'ha == wPos) begin
            mem_10 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'ha == _T_308) begin
                mem_10 <= _GEN_31;
              end else begin
                if (6'ha == _T_303) begin
                  mem_10 <= _GEN_30;
                end else begin
                  if (6'ha == _T_298) begin
                    mem_10 <= _GEN_29;
                  end else begin
                    if (6'ha == _T_293) begin
                      mem_10 <= _GEN_28;
                    end else begin
                      if (6'ha == _T_288) begin
                        mem_10 <= _GEN_27;
                      end else begin
                        if (6'ha == _T_283) begin
                          mem_10 <= _GEN_26;
                        end else begin
                          if (6'ha == _T_278) begin
                            mem_10 <= _GEN_25;
                          end else begin
                            if (6'ha == _T_273) begin
                              mem_10 <= _GEN_24;
                            end else begin
                              if (6'ha == _T_268) begin
                                mem_10 <= _GEN_23;
                              end else begin
                                if (6'ha == _T_263) begin
                                  mem_10 <= _GEN_22;
                                end else begin
                                  if (6'ha == _T_258) begin
                                    mem_10 <= _GEN_21;
                                  end else begin
                                    if (6'ha == _T_253) begin
                                      mem_10 <= _GEN_20;
                                    end else begin
                                      if (6'ha == _T_248) begin
                                        mem_10 <= _GEN_19;
                                      end else begin
                                        if (6'ha == _T_243) begin
                                          mem_10 <= _GEN_18;
                                        end else begin
                                          if (6'ha == _T_238) begin
                                            mem_10 <= _GEN_17;
                                          end else begin
                                            if (6'ha == _T_233) begin
                                              mem_10 <= _GEN_16;
                                            end else begin
                                              if (6'ha == _T_228) begin
                                                mem_10 <= _GEN_15;
                                              end else begin
                                                if (6'ha == _T_223) begin
                                                  mem_10 <= _GEN_14;
                                                end else begin
                                                  if (6'ha == _T_218) begin
                                                    mem_10 <= _GEN_13;
                                                  end else begin
                                                    if (6'ha == _T_213) begin
                                                      mem_10 <= _GEN_12;
                                                    end else begin
                                                      if (6'ha == _T_208) begin
                                                        mem_10 <= _GEN_11;
                                                      end else begin
                                                        if (6'ha == _T_203) begin
                                                          mem_10 <= _GEN_10;
                                                        end else begin
                                                          if (6'ha == _T_198) begin
                                                            mem_10 <= _GEN_9;
                                                          end else begin
                                                            if (6'ha == _T_193) begin
                                                              mem_10 <= _GEN_8;
                                                            end else begin
                                                              if (6'ha == _T_188) begin
                                                                mem_10 <= _GEN_7;
                                                              end else begin
                                                                if (6'ha == _T_183) begin
                                                                  mem_10 <= _GEN_6;
                                                                end else begin
                                                                  if (6'ha == _T_178) begin
                                                                    mem_10 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'ha == _T_173) begin
                                                                      mem_10 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'ha == _T_168) begin
                                                                        mem_10 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'ha == _T_163) begin
                                                                          mem_10 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'ha == _T_158) begin
                                                                            mem_10 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'ha == _T_153) begin
                                                                              mem_10 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'ha == _T_308) begin
              mem_10 <= _GEN_31;
            end else begin
              if (6'ha == _T_303) begin
                mem_10 <= _GEN_30;
              end else begin
                if (6'ha == _T_298) begin
                  mem_10 <= _GEN_29;
                end else begin
                  if (6'ha == _T_293) begin
                    mem_10 <= _GEN_28;
                  end else begin
                    if (6'ha == _T_288) begin
                      mem_10 <= _GEN_27;
                    end else begin
                      if (6'ha == _T_283) begin
                        mem_10 <= _GEN_26;
                      end else begin
                        if (6'ha == _T_278) begin
                          mem_10 <= _GEN_25;
                        end else begin
                          if (6'ha == _T_273) begin
                            mem_10 <= _GEN_24;
                          end else begin
                            if (6'ha == _T_268) begin
                              mem_10 <= _GEN_23;
                            end else begin
                              if (6'ha == _T_263) begin
                                mem_10 <= _GEN_22;
                              end else begin
                                if (6'ha == _T_258) begin
                                  mem_10 <= _GEN_21;
                                end else begin
                                  if (6'ha == _T_253) begin
                                    mem_10 <= _GEN_20;
                                  end else begin
                                    if (6'ha == _T_248) begin
                                      mem_10 <= _GEN_19;
                                    end else begin
                                      if (6'ha == _T_243) begin
                                        mem_10 <= _GEN_18;
                                      end else begin
                                        if (6'ha == _T_238) begin
                                          mem_10 <= _GEN_17;
                                        end else begin
                                          if (6'ha == _T_233) begin
                                            mem_10 <= _GEN_16;
                                          end else begin
                                            if (6'ha == _T_228) begin
                                              mem_10 <= _GEN_15;
                                            end else begin
                                              if (6'ha == _T_223) begin
                                                mem_10 <= _GEN_14;
                                              end else begin
                                                if (6'ha == _T_218) begin
                                                  mem_10 <= _GEN_13;
                                                end else begin
                                                  if (6'ha == _T_213) begin
                                                    mem_10 <= _GEN_12;
                                                  end else begin
                                                    if (6'ha == _T_208) begin
                                                      mem_10 <= _GEN_11;
                                                    end else begin
                                                      if (6'ha == _T_203) begin
                                                        mem_10 <= _GEN_10;
                                                      end else begin
                                                        if (6'ha == _T_198) begin
                                                          mem_10 <= _GEN_9;
                                                        end else begin
                                                          if (6'ha == _T_193) begin
                                                            mem_10 <= _GEN_8;
                                                          end else begin
                                                            if (6'ha == _T_188) begin
                                                              mem_10 <= _GEN_7;
                                                            end else begin
                                                              if (6'ha == _T_183) begin
                                                                mem_10 <= _GEN_6;
                                                              end else begin
                                                                if (6'ha == _T_178) begin
                                                                  mem_10 <= _GEN_5;
                                                                end else begin
                                                                  if (6'ha == _T_173) begin
                                                                    mem_10 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'ha == _T_168) begin
                                                                      mem_10 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'ha == _T_163) begin
                                                                        mem_10 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'ha == _T_158) begin
                                                                          mem_10 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'ha == _T_153) begin
                                                                            mem_10 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'ha == _T_308) begin
            mem_10 <= _GEN_31;
          end else begin
            if (6'ha == _T_303) begin
              mem_10 <= _GEN_30;
            end else begin
              if (6'ha == _T_298) begin
                mem_10 <= _GEN_29;
              end else begin
                if (6'ha == _T_293) begin
                  mem_10 <= _GEN_28;
                end else begin
                  if (6'ha == _T_288) begin
                    mem_10 <= _GEN_27;
                  end else begin
                    if (6'ha == _T_283) begin
                      mem_10 <= _GEN_26;
                    end else begin
                      if (6'ha == _T_278) begin
                        mem_10 <= _GEN_25;
                      end else begin
                        if (6'ha == _T_273) begin
                          mem_10 <= _GEN_24;
                        end else begin
                          if (6'ha == _T_268) begin
                            mem_10 <= _GEN_23;
                          end else begin
                            if (6'ha == _T_263) begin
                              mem_10 <= _GEN_22;
                            end else begin
                              if (6'ha == _T_258) begin
                                mem_10 <= _GEN_21;
                              end else begin
                                if (6'ha == _T_253) begin
                                  mem_10 <= _GEN_20;
                                end else begin
                                  if (6'ha == _T_248) begin
                                    mem_10 <= _GEN_19;
                                  end else begin
                                    if (6'ha == _T_243) begin
                                      mem_10 <= _GEN_18;
                                    end else begin
                                      if (6'ha == _T_238) begin
                                        mem_10 <= _GEN_17;
                                      end else begin
                                        if (6'ha == _T_233) begin
                                          mem_10 <= _GEN_16;
                                        end else begin
                                          if (6'ha == _T_228) begin
                                            mem_10 <= _GEN_15;
                                          end else begin
                                            if (6'ha == _T_223) begin
                                              mem_10 <= _GEN_14;
                                            end else begin
                                              if (6'ha == _T_218) begin
                                                mem_10 <= _GEN_13;
                                              end else begin
                                                if (6'ha == _T_213) begin
                                                  mem_10 <= _GEN_12;
                                                end else begin
                                                  if (6'ha == _T_208) begin
                                                    mem_10 <= _GEN_11;
                                                  end else begin
                                                    if (6'ha == _T_203) begin
                                                      mem_10 <= _GEN_10;
                                                    end else begin
                                                      if (6'ha == _T_198) begin
                                                        mem_10 <= _GEN_9;
                                                      end else begin
                                                        if (6'ha == _T_193) begin
                                                          mem_10 <= _GEN_8;
                                                        end else begin
                                                          if (6'ha == _T_188) begin
                                                            mem_10 <= _GEN_7;
                                                          end else begin
                                                            if (6'ha == _T_183) begin
                                                              mem_10 <= _GEN_6;
                                                            end else begin
                                                              if (6'ha == _T_178) begin
                                                                mem_10 <= _GEN_5;
                                                              end else begin
                                                                if (6'ha == _T_173) begin
                                                                  mem_10 <= _GEN_4;
                                                                end else begin
                                                                  if (6'ha == _T_168) begin
                                                                    mem_10 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'ha == _T_163) begin
                                                                      mem_10 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'ha == _T_158) begin
                                                                        mem_10 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'ha == _T_153) begin
                                                                          mem_10 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'ha == _T_308) begin
          mem_10 <= _GEN_31;
        end else begin
          if (6'ha == _T_303) begin
            mem_10 <= _GEN_30;
          end else begin
            if (6'ha == _T_298) begin
              mem_10 <= _GEN_29;
            end else begin
              if (6'ha == _T_293) begin
                mem_10 <= _GEN_28;
              end else begin
                if (6'ha == _T_288) begin
                  mem_10 <= _GEN_27;
                end else begin
                  if (6'ha == _T_283) begin
                    mem_10 <= _GEN_26;
                  end else begin
                    if (6'ha == _T_278) begin
                      mem_10 <= _GEN_25;
                    end else begin
                      if (6'ha == _T_273) begin
                        mem_10 <= _GEN_24;
                      end else begin
                        if (6'ha == _T_268) begin
                          mem_10 <= _GEN_23;
                        end else begin
                          if (6'ha == _T_263) begin
                            mem_10 <= _GEN_22;
                          end else begin
                            if (6'ha == _T_258) begin
                              mem_10 <= _GEN_21;
                            end else begin
                              if (6'ha == _T_253) begin
                                mem_10 <= _GEN_20;
                              end else begin
                                if (6'ha == _T_248) begin
                                  mem_10 <= _GEN_19;
                                end else begin
                                  if (6'ha == _T_243) begin
                                    mem_10 <= _GEN_18;
                                  end else begin
                                    if (6'ha == _T_238) begin
                                      mem_10 <= _GEN_17;
                                    end else begin
                                      if (6'ha == _T_233) begin
                                        mem_10 <= _GEN_16;
                                      end else begin
                                        if (6'ha == _T_228) begin
                                          mem_10 <= _GEN_15;
                                        end else begin
                                          if (6'ha == _T_223) begin
                                            mem_10 <= _GEN_14;
                                          end else begin
                                            if (6'ha == _T_218) begin
                                              mem_10 <= _GEN_13;
                                            end else begin
                                              if (6'ha == _T_213) begin
                                                mem_10 <= _GEN_12;
                                              end else begin
                                                if (6'ha == _T_208) begin
                                                  mem_10 <= _GEN_11;
                                                end else begin
                                                  if (6'ha == _T_203) begin
                                                    mem_10 <= _GEN_10;
                                                  end else begin
                                                    if (6'ha == _T_198) begin
                                                      mem_10 <= _GEN_9;
                                                    end else begin
                                                      if (6'ha == _T_193) begin
                                                        mem_10 <= _GEN_8;
                                                      end else begin
                                                        if (6'ha == _T_188) begin
                                                          mem_10 <= _GEN_7;
                                                        end else begin
                                                          if (6'ha == _T_183) begin
                                                            mem_10 <= _GEN_6;
                                                          end else begin
                                                            if (6'ha == _T_178) begin
                                                              mem_10 <= _GEN_5;
                                                            end else begin
                                                              if (6'ha == _T_173) begin
                                                                mem_10 <= _GEN_4;
                                                              end else begin
                                                                if (6'ha == _T_168) begin
                                                                  mem_10 <= _GEN_3;
                                                                end else begin
                                                                  if (6'ha == _T_163) begin
                                                                    mem_10 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'ha == _T_158) begin
                                                                      mem_10 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'ha == _T_153) begin
                                                                        mem_10 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'hb == wPos) begin
            mem_11 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'hb == _T_308) begin
                mem_11 <= _GEN_31;
              end else begin
                if (6'hb == _T_303) begin
                  mem_11 <= _GEN_30;
                end else begin
                  if (6'hb == _T_298) begin
                    mem_11 <= _GEN_29;
                  end else begin
                    if (6'hb == _T_293) begin
                      mem_11 <= _GEN_28;
                    end else begin
                      if (6'hb == _T_288) begin
                        mem_11 <= _GEN_27;
                      end else begin
                        if (6'hb == _T_283) begin
                          mem_11 <= _GEN_26;
                        end else begin
                          if (6'hb == _T_278) begin
                            mem_11 <= _GEN_25;
                          end else begin
                            if (6'hb == _T_273) begin
                              mem_11 <= _GEN_24;
                            end else begin
                              if (6'hb == _T_268) begin
                                mem_11 <= _GEN_23;
                              end else begin
                                if (6'hb == _T_263) begin
                                  mem_11 <= _GEN_22;
                                end else begin
                                  if (6'hb == _T_258) begin
                                    mem_11 <= _GEN_21;
                                  end else begin
                                    if (6'hb == _T_253) begin
                                      mem_11 <= _GEN_20;
                                    end else begin
                                      if (6'hb == _T_248) begin
                                        mem_11 <= _GEN_19;
                                      end else begin
                                        if (6'hb == _T_243) begin
                                          mem_11 <= _GEN_18;
                                        end else begin
                                          if (6'hb == _T_238) begin
                                            mem_11 <= _GEN_17;
                                          end else begin
                                            if (6'hb == _T_233) begin
                                              mem_11 <= _GEN_16;
                                            end else begin
                                              if (6'hb == _T_228) begin
                                                mem_11 <= _GEN_15;
                                              end else begin
                                                if (6'hb == _T_223) begin
                                                  mem_11 <= _GEN_14;
                                                end else begin
                                                  if (6'hb == _T_218) begin
                                                    mem_11 <= _GEN_13;
                                                  end else begin
                                                    if (6'hb == _T_213) begin
                                                      mem_11 <= _GEN_12;
                                                    end else begin
                                                      if (6'hb == _T_208) begin
                                                        mem_11 <= _GEN_11;
                                                      end else begin
                                                        if (6'hb == _T_203) begin
                                                          mem_11 <= _GEN_10;
                                                        end else begin
                                                          if (6'hb == _T_198) begin
                                                            mem_11 <= _GEN_9;
                                                          end else begin
                                                            if (6'hb == _T_193) begin
                                                              mem_11 <= _GEN_8;
                                                            end else begin
                                                              if (6'hb == _T_188) begin
                                                                mem_11 <= _GEN_7;
                                                              end else begin
                                                                if (6'hb == _T_183) begin
                                                                  mem_11 <= _GEN_6;
                                                                end else begin
                                                                  if (6'hb == _T_178) begin
                                                                    mem_11 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'hb == _T_173) begin
                                                                      mem_11 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'hb == _T_168) begin
                                                                        mem_11 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'hb == _T_163) begin
                                                                          mem_11 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'hb == _T_158) begin
                                                                            mem_11 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'hb == _T_153) begin
                                                                              mem_11 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'hb == _T_308) begin
              mem_11 <= _GEN_31;
            end else begin
              if (6'hb == _T_303) begin
                mem_11 <= _GEN_30;
              end else begin
                if (6'hb == _T_298) begin
                  mem_11 <= _GEN_29;
                end else begin
                  if (6'hb == _T_293) begin
                    mem_11 <= _GEN_28;
                  end else begin
                    if (6'hb == _T_288) begin
                      mem_11 <= _GEN_27;
                    end else begin
                      if (6'hb == _T_283) begin
                        mem_11 <= _GEN_26;
                      end else begin
                        if (6'hb == _T_278) begin
                          mem_11 <= _GEN_25;
                        end else begin
                          if (6'hb == _T_273) begin
                            mem_11 <= _GEN_24;
                          end else begin
                            if (6'hb == _T_268) begin
                              mem_11 <= _GEN_23;
                            end else begin
                              if (6'hb == _T_263) begin
                                mem_11 <= _GEN_22;
                              end else begin
                                if (6'hb == _T_258) begin
                                  mem_11 <= _GEN_21;
                                end else begin
                                  if (6'hb == _T_253) begin
                                    mem_11 <= _GEN_20;
                                  end else begin
                                    if (6'hb == _T_248) begin
                                      mem_11 <= _GEN_19;
                                    end else begin
                                      if (6'hb == _T_243) begin
                                        mem_11 <= _GEN_18;
                                      end else begin
                                        if (6'hb == _T_238) begin
                                          mem_11 <= _GEN_17;
                                        end else begin
                                          if (6'hb == _T_233) begin
                                            mem_11 <= _GEN_16;
                                          end else begin
                                            if (6'hb == _T_228) begin
                                              mem_11 <= _GEN_15;
                                            end else begin
                                              if (6'hb == _T_223) begin
                                                mem_11 <= _GEN_14;
                                              end else begin
                                                if (6'hb == _T_218) begin
                                                  mem_11 <= _GEN_13;
                                                end else begin
                                                  if (6'hb == _T_213) begin
                                                    mem_11 <= _GEN_12;
                                                  end else begin
                                                    if (6'hb == _T_208) begin
                                                      mem_11 <= _GEN_11;
                                                    end else begin
                                                      if (6'hb == _T_203) begin
                                                        mem_11 <= _GEN_10;
                                                      end else begin
                                                        if (6'hb == _T_198) begin
                                                          mem_11 <= _GEN_9;
                                                        end else begin
                                                          if (6'hb == _T_193) begin
                                                            mem_11 <= _GEN_8;
                                                          end else begin
                                                            if (6'hb == _T_188) begin
                                                              mem_11 <= _GEN_7;
                                                            end else begin
                                                              if (6'hb == _T_183) begin
                                                                mem_11 <= _GEN_6;
                                                              end else begin
                                                                if (6'hb == _T_178) begin
                                                                  mem_11 <= _GEN_5;
                                                                end else begin
                                                                  if (6'hb == _T_173) begin
                                                                    mem_11 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'hb == _T_168) begin
                                                                      mem_11 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'hb == _T_163) begin
                                                                        mem_11 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'hb == _T_158) begin
                                                                          mem_11 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'hb == _T_153) begin
                                                                            mem_11 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'hb == _T_308) begin
            mem_11 <= _GEN_31;
          end else begin
            if (6'hb == _T_303) begin
              mem_11 <= _GEN_30;
            end else begin
              if (6'hb == _T_298) begin
                mem_11 <= _GEN_29;
              end else begin
                if (6'hb == _T_293) begin
                  mem_11 <= _GEN_28;
                end else begin
                  if (6'hb == _T_288) begin
                    mem_11 <= _GEN_27;
                  end else begin
                    if (6'hb == _T_283) begin
                      mem_11 <= _GEN_26;
                    end else begin
                      if (6'hb == _T_278) begin
                        mem_11 <= _GEN_25;
                      end else begin
                        if (6'hb == _T_273) begin
                          mem_11 <= _GEN_24;
                        end else begin
                          if (6'hb == _T_268) begin
                            mem_11 <= _GEN_23;
                          end else begin
                            if (6'hb == _T_263) begin
                              mem_11 <= _GEN_22;
                            end else begin
                              if (6'hb == _T_258) begin
                                mem_11 <= _GEN_21;
                              end else begin
                                if (6'hb == _T_253) begin
                                  mem_11 <= _GEN_20;
                                end else begin
                                  if (6'hb == _T_248) begin
                                    mem_11 <= _GEN_19;
                                  end else begin
                                    if (6'hb == _T_243) begin
                                      mem_11 <= _GEN_18;
                                    end else begin
                                      if (6'hb == _T_238) begin
                                        mem_11 <= _GEN_17;
                                      end else begin
                                        if (6'hb == _T_233) begin
                                          mem_11 <= _GEN_16;
                                        end else begin
                                          if (6'hb == _T_228) begin
                                            mem_11 <= _GEN_15;
                                          end else begin
                                            if (6'hb == _T_223) begin
                                              mem_11 <= _GEN_14;
                                            end else begin
                                              if (6'hb == _T_218) begin
                                                mem_11 <= _GEN_13;
                                              end else begin
                                                if (6'hb == _T_213) begin
                                                  mem_11 <= _GEN_12;
                                                end else begin
                                                  if (6'hb == _T_208) begin
                                                    mem_11 <= _GEN_11;
                                                  end else begin
                                                    if (6'hb == _T_203) begin
                                                      mem_11 <= _GEN_10;
                                                    end else begin
                                                      if (6'hb == _T_198) begin
                                                        mem_11 <= _GEN_9;
                                                      end else begin
                                                        if (6'hb == _T_193) begin
                                                          mem_11 <= _GEN_8;
                                                        end else begin
                                                          if (6'hb == _T_188) begin
                                                            mem_11 <= _GEN_7;
                                                          end else begin
                                                            if (6'hb == _T_183) begin
                                                              mem_11 <= _GEN_6;
                                                            end else begin
                                                              if (6'hb == _T_178) begin
                                                                mem_11 <= _GEN_5;
                                                              end else begin
                                                                if (6'hb == _T_173) begin
                                                                  mem_11 <= _GEN_4;
                                                                end else begin
                                                                  if (6'hb == _T_168) begin
                                                                    mem_11 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'hb == _T_163) begin
                                                                      mem_11 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'hb == _T_158) begin
                                                                        mem_11 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'hb == _T_153) begin
                                                                          mem_11 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'hb == _T_308) begin
          mem_11 <= _GEN_31;
        end else begin
          if (6'hb == _T_303) begin
            mem_11 <= _GEN_30;
          end else begin
            if (6'hb == _T_298) begin
              mem_11 <= _GEN_29;
            end else begin
              if (6'hb == _T_293) begin
                mem_11 <= _GEN_28;
              end else begin
                if (6'hb == _T_288) begin
                  mem_11 <= _GEN_27;
                end else begin
                  if (6'hb == _T_283) begin
                    mem_11 <= _GEN_26;
                  end else begin
                    if (6'hb == _T_278) begin
                      mem_11 <= _GEN_25;
                    end else begin
                      if (6'hb == _T_273) begin
                        mem_11 <= _GEN_24;
                      end else begin
                        if (6'hb == _T_268) begin
                          mem_11 <= _GEN_23;
                        end else begin
                          if (6'hb == _T_263) begin
                            mem_11 <= _GEN_22;
                          end else begin
                            if (6'hb == _T_258) begin
                              mem_11 <= _GEN_21;
                            end else begin
                              if (6'hb == _T_253) begin
                                mem_11 <= _GEN_20;
                              end else begin
                                if (6'hb == _T_248) begin
                                  mem_11 <= _GEN_19;
                                end else begin
                                  if (6'hb == _T_243) begin
                                    mem_11 <= _GEN_18;
                                  end else begin
                                    if (6'hb == _T_238) begin
                                      mem_11 <= _GEN_17;
                                    end else begin
                                      if (6'hb == _T_233) begin
                                        mem_11 <= _GEN_16;
                                      end else begin
                                        if (6'hb == _T_228) begin
                                          mem_11 <= _GEN_15;
                                        end else begin
                                          if (6'hb == _T_223) begin
                                            mem_11 <= _GEN_14;
                                          end else begin
                                            if (6'hb == _T_218) begin
                                              mem_11 <= _GEN_13;
                                            end else begin
                                              if (6'hb == _T_213) begin
                                                mem_11 <= _GEN_12;
                                              end else begin
                                                if (6'hb == _T_208) begin
                                                  mem_11 <= _GEN_11;
                                                end else begin
                                                  if (6'hb == _T_203) begin
                                                    mem_11 <= _GEN_10;
                                                  end else begin
                                                    if (6'hb == _T_198) begin
                                                      mem_11 <= _GEN_9;
                                                    end else begin
                                                      if (6'hb == _T_193) begin
                                                        mem_11 <= _GEN_8;
                                                      end else begin
                                                        if (6'hb == _T_188) begin
                                                          mem_11 <= _GEN_7;
                                                        end else begin
                                                          if (6'hb == _T_183) begin
                                                            mem_11 <= _GEN_6;
                                                          end else begin
                                                            if (6'hb == _T_178) begin
                                                              mem_11 <= _GEN_5;
                                                            end else begin
                                                              if (6'hb == _T_173) begin
                                                                mem_11 <= _GEN_4;
                                                              end else begin
                                                                if (6'hb == _T_168) begin
                                                                  mem_11 <= _GEN_3;
                                                                end else begin
                                                                  if (6'hb == _T_163) begin
                                                                    mem_11 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'hb == _T_158) begin
                                                                      mem_11 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'hb == _T_153) begin
                                                                        mem_11 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'hc == wPos) begin
            mem_12 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'hc == _T_308) begin
                mem_12 <= _GEN_31;
              end else begin
                if (6'hc == _T_303) begin
                  mem_12 <= _GEN_30;
                end else begin
                  if (6'hc == _T_298) begin
                    mem_12 <= _GEN_29;
                  end else begin
                    if (6'hc == _T_293) begin
                      mem_12 <= _GEN_28;
                    end else begin
                      if (6'hc == _T_288) begin
                        mem_12 <= _GEN_27;
                      end else begin
                        if (6'hc == _T_283) begin
                          mem_12 <= _GEN_26;
                        end else begin
                          if (6'hc == _T_278) begin
                            mem_12 <= _GEN_25;
                          end else begin
                            if (6'hc == _T_273) begin
                              mem_12 <= _GEN_24;
                            end else begin
                              if (6'hc == _T_268) begin
                                mem_12 <= _GEN_23;
                              end else begin
                                if (6'hc == _T_263) begin
                                  mem_12 <= _GEN_22;
                                end else begin
                                  if (6'hc == _T_258) begin
                                    mem_12 <= _GEN_21;
                                  end else begin
                                    if (6'hc == _T_253) begin
                                      mem_12 <= _GEN_20;
                                    end else begin
                                      if (6'hc == _T_248) begin
                                        mem_12 <= _GEN_19;
                                      end else begin
                                        if (6'hc == _T_243) begin
                                          mem_12 <= _GEN_18;
                                        end else begin
                                          if (6'hc == _T_238) begin
                                            mem_12 <= _GEN_17;
                                          end else begin
                                            if (6'hc == _T_233) begin
                                              mem_12 <= _GEN_16;
                                            end else begin
                                              if (6'hc == _T_228) begin
                                                mem_12 <= _GEN_15;
                                              end else begin
                                                if (6'hc == _T_223) begin
                                                  mem_12 <= _GEN_14;
                                                end else begin
                                                  if (6'hc == _T_218) begin
                                                    mem_12 <= _GEN_13;
                                                  end else begin
                                                    if (6'hc == _T_213) begin
                                                      mem_12 <= _GEN_12;
                                                    end else begin
                                                      if (6'hc == _T_208) begin
                                                        mem_12 <= _GEN_11;
                                                      end else begin
                                                        if (6'hc == _T_203) begin
                                                          mem_12 <= _GEN_10;
                                                        end else begin
                                                          if (6'hc == _T_198) begin
                                                            mem_12 <= _GEN_9;
                                                          end else begin
                                                            if (6'hc == _T_193) begin
                                                              mem_12 <= _GEN_8;
                                                            end else begin
                                                              if (6'hc == _T_188) begin
                                                                mem_12 <= _GEN_7;
                                                              end else begin
                                                                if (6'hc == _T_183) begin
                                                                  mem_12 <= _GEN_6;
                                                                end else begin
                                                                  if (6'hc == _T_178) begin
                                                                    mem_12 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'hc == _T_173) begin
                                                                      mem_12 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'hc == _T_168) begin
                                                                        mem_12 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'hc == _T_163) begin
                                                                          mem_12 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'hc == _T_158) begin
                                                                            mem_12 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'hc == _T_153) begin
                                                                              mem_12 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'hc == _T_308) begin
              mem_12 <= _GEN_31;
            end else begin
              if (6'hc == _T_303) begin
                mem_12 <= _GEN_30;
              end else begin
                if (6'hc == _T_298) begin
                  mem_12 <= _GEN_29;
                end else begin
                  if (6'hc == _T_293) begin
                    mem_12 <= _GEN_28;
                  end else begin
                    if (6'hc == _T_288) begin
                      mem_12 <= _GEN_27;
                    end else begin
                      if (6'hc == _T_283) begin
                        mem_12 <= _GEN_26;
                      end else begin
                        if (6'hc == _T_278) begin
                          mem_12 <= _GEN_25;
                        end else begin
                          if (6'hc == _T_273) begin
                            mem_12 <= _GEN_24;
                          end else begin
                            if (6'hc == _T_268) begin
                              mem_12 <= _GEN_23;
                            end else begin
                              if (6'hc == _T_263) begin
                                mem_12 <= _GEN_22;
                              end else begin
                                if (6'hc == _T_258) begin
                                  mem_12 <= _GEN_21;
                                end else begin
                                  if (6'hc == _T_253) begin
                                    mem_12 <= _GEN_20;
                                  end else begin
                                    if (6'hc == _T_248) begin
                                      mem_12 <= _GEN_19;
                                    end else begin
                                      if (6'hc == _T_243) begin
                                        mem_12 <= _GEN_18;
                                      end else begin
                                        if (6'hc == _T_238) begin
                                          mem_12 <= _GEN_17;
                                        end else begin
                                          if (6'hc == _T_233) begin
                                            mem_12 <= _GEN_16;
                                          end else begin
                                            if (6'hc == _T_228) begin
                                              mem_12 <= _GEN_15;
                                            end else begin
                                              if (6'hc == _T_223) begin
                                                mem_12 <= _GEN_14;
                                              end else begin
                                                if (6'hc == _T_218) begin
                                                  mem_12 <= _GEN_13;
                                                end else begin
                                                  if (6'hc == _T_213) begin
                                                    mem_12 <= _GEN_12;
                                                  end else begin
                                                    if (6'hc == _T_208) begin
                                                      mem_12 <= _GEN_11;
                                                    end else begin
                                                      if (6'hc == _T_203) begin
                                                        mem_12 <= _GEN_10;
                                                      end else begin
                                                        if (6'hc == _T_198) begin
                                                          mem_12 <= _GEN_9;
                                                        end else begin
                                                          if (6'hc == _T_193) begin
                                                            mem_12 <= _GEN_8;
                                                          end else begin
                                                            if (6'hc == _T_188) begin
                                                              mem_12 <= _GEN_7;
                                                            end else begin
                                                              if (6'hc == _T_183) begin
                                                                mem_12 <= _GEN_6;
                                                              end else begin
                                                                if (6'hc == _T_178) begin
                                                                  mem_12 <= _GEN_5;
                                                                end else begin
                                                                  if (6'hc == _T_173) begin
                                                                    mem_12 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'hc == _T_168) begin
                                                                      mem_12 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'hc == _T_163) begin
                                                                        mem_12 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'hc == _T_158) begin
                                                                          mem_12 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'hc == _T_153) begin
                                                                            mem_12 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'hc == _T_308) begin
            mem_12 <= _GEN_31;
          end else begin
            if (6'hc == _T_303) begin
              mem_12 <= _GEN_30;
            end else begin
              if (6'hc == _T_298) begin
                mem_12 <= _GEN_29;
              end else begin
                if (6'hc == _T_293) begin
                  mem_12 <= _GEN_28;
                end else begin
                  if (6'hc == _T_288) begin
                    mem_12 <= _GEN_27;
                  end else begin
                    if (6'hc == _T_283) begin
                      mem_12 <= _GEN_26;
                    end else begin
                      if (6'hc == _T_278) begin
                        mem_12 <= _GEN_25;
                      end else begin
                        if (6'hc == _T_273) begin
                          mem_12 <= _GEN_24;
                        end else begin
                          if (6'hc == _T_268) begin
                            mem_12 <= _GEN_23;
                          end else begin
                            if (6'hc == _T_263) begin
                              mem_12 <= _GEN_22;
                            end else begin
                              if (6'hc == _T_258) begin
                                mem_12 <= _GEN_21;
                              end else begin
                                if (6'hc == _T_253) begin
                                  mem_12 <= _GEN_20;
                                end else begin
                                  if (6'hc == _T_248) begin
                                    mem_12 <= _GEN_19;
                                  end else begin
                                    if (6'hc == _T_243) begin
                                      mem_12 <= _GEN_18;
                                    end else begin
                                      if (6'hc == _T_238) begin
                                        mem_12 <= _GEN_17;
                                      end else begin
                                        if (6'hc == _T_233) begin
                                          mem_12 <= _GEN_16;
                                        end else begin
                                          if (6'hc == _T_228) begin
                                            mem_12 <= _GEN_15;
                                          end else begin
                                            if (6'hc == _T_223) begin
                                              mem_12 <= _GEN_14;
                                            end else begin
                                              if (6'hc == _T_218) begin
                                                mem_12 <= _GEN_13;
                                              end else begin
                                                if (6'hc == _T_213) begin
                                                  mem_12 <= _GEN_12;
                                                end else begin
                                                  if (6'hc == _T_208) begin
                                                    mem_12 <= _GEN_11;
                                                  end else begin
                                                    if (6'hc == _T_203) begin
                                                      mem_12 <= _GEN_10;
                                                    end else begin
                                                      if (6'hc == _T_198) begin
                                                        mem_12 <= _GEN_9;
                                                      end else begin
                                                        if (6'hc == _T_193) begin
                                                          mem_12 <= _GEN_8;
                                                        end else begin
                                                          if (6'hc == _T_188) begin
                                                            mem_12 <= _GEN_7;
                                                          end else begin
                                                            if (6'hc == _T_183) begin
                                                              mem_12 <= _GEN_6;
                                                            end else begin
                                                              if (6'hc == _T_178) begin
                                                                mem_12 <= _GEN_5;
                                                              end else begin
                                                                if (6'hc == _T_173) begin
                                                                  mem_12 <= _GEN_4;
                                                                end else begin
                                                                  if (6'hc == _T_168) begin
                                                                    mem_12 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'hc == _T_163) begin
                                                                      mem_12 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'hc == _T_158) begin
                                                                        mem_12 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'hc == _T_153) begin
                                                                          mem_12 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'hc == _T_308) begin
          mem_12 <= _GEN_31;
        end else begin
          if (6'hc == _T_303) begin
            mem_12 <= _GEN_30;
          end else begin
            if (6'hc == _T_298) begin
              mem_12 <= _GEN_29;
            end else begin
              if (6'hc == _T_293) begin
                mem_12 <= _GEN_28;
              end else begin
                if (6'hc == _T_288) begin
                  mem_12 <= _GEN_27;
                end else begin
                  if (6'hc == _T_283) begin
                    mem_12 <= _GEN_26;
                  end else begin
                    if (6'hc == _T_278) begin
                      mem_12 <= _GEN_25;
                    end else begin
                      if (6'hc == _T_273) begin
                        mem_12 <= _GEN_24;
                      end else begin
                        if (6'hc == _T_268) begin
                          mem_12 <= _GEN_23;
                        end else begin
                          if (6'hc == _T_263) begin
                            mem_12 <= _GEN_22;
                          end else begin
                            if (6'hc == _T_258) begin
                              mem_12 <= _GEN_21;
                            end else begin
                              if (6'hc == _T_253) begin
                                mem_12 <= _GEN_20;
                              end else begin
                                if (6'hc == _T_248) begin
                                  mem_12 <= _GEN_19;
                                end else begin
                                  if (6'hc == _T_243) begin
                                    mem_12 <= _GEN_18;
                                  end else begin
                                    if (6'hc == _T_238) begin
                                      mem_12 <= _GEN_17;
                                    end else begin
                                      if (6'hc == _T_233) begin
                                        mem_12 <= _GEN_16;
                                      end else begin
                                        if (6'hc == _T_228) begin
                                          mem_12 <= _GEN_15;
                                        end else begin
                                          if (6'hc == _T_223) begin
                                            mem_12 <= _GEN_14;
                                          end else begin
                                            if (6'hc == _T_218) begin
                                              mem_12 <= _GEN_13;
                                            end else begin
                                              if (6'hc == _T_213) begin
                                                mem_12 <= _GEN_12;
                                              end else begin
                                                if (6'hc == _T_208) begin
                                                  mem_12 <= _GEN_11;
                                                end else begin
                                                  if (6'hc == _T_203) begin
                                                    mem_12 <= _GEN_10;
                                                  end else begin
                                                    if (6'hc == _T_198) begin
                                                      mem_12 <= _GEN_9;
                                                    end else begin
                                                      if (6'hc == _T_193) begin
                                                        mem_12 <= _GEN_8;
                                                      end else begin
                                                        if (6'hc == _T_188) begin
                                                          mem_12 <= _GEN_7;
                                                        end else begin
                                                          if (6'hc == _T_183) begin
                                                            mem_12 <= _GEN_6;
                                                          end else begin
                                                            if (6'hc == _T_178) begin
                                                              mem_12 <= _GEN_5;
                                                            end else begin
                                                              if (6'hc == _T_173) begin
                                                                mem_12 <= _GEN_4;
                                                              end else begin
                                                                if (6'hc == _T_168) begin
                                                                  mem_12 <= _GEN_3;
                                                                end else begin
                                                                  if (6'hc == _T_163) begin
                                                                    mem_12 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'hc == _T_158) begin
                                                                      mem_12 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'hc == _T_153) begin
                                                                        mem_12 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'hd == wPos) begin
            mem_13 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'hd == _T_308) begin
                mem_13 <= _GEN_31;
              end else begin
                if (6'hd == _T_303) begin
                  mem_13 <= _GEN_30;
                end else begin
                  if (6'hd == _T_298) begin
                    mem_13 <= _GEN_29;
                  end else begin
                    if (6'hd == _T_293) begin
                      mem_13 <= _GEN_28;
                    end else begin
                      if (6'hd == _T_288) begin
                        mem_13 <= _GEN_27;
                      end else begin
                        if (6'hd == _T_283) begin
                          mem_13 <= _GEN_26;
                        end else begin
                          if (6'hd == _T_278) begin
                            mem_13 <= _GEN_25;
                          end else begin
                            if (6'hd == _T_273) begin
                              mem_13 <= _GEN_24;
                            end else begin
                              if (6'hd == _T_268) begin
                                mem_13 <= _GEN_23;
                              end else begin
                                if (6'hd == _T_263) begin
                                  mem_13 <= _GEN_22;
                                end else begin
                                  if (6'hd == _T_258) begin
                                    mem_13 <= _GEN_21;
                                  end else begin
                                    if (6'hd == _T_253) begin
                                      mem_13 <= _GEN_20;
                                    end else begin
                                      if (6'hd == _T_248) begin
                                        mem_13 <= _GEN_19;
                                      end else begin
                                        if (6'hd == _T_243) begin
                                          mem_13 <= _GEN_18;
                                        end else begin
                                          if (6'hd == _T_238) begin
                                            mem_13 <= _GEN_17;
                                          end else begin
                                            if (6'hd == _T_233) begin
                                              mem_13 <= _GEN_16;
                                            end else begin
                                              if (6'hd == _T_228) begin
                                                mem_13 <= _GEN_15;
                                              end else begin
                                                if (6'hd == _T_223) begin
                                                  mem_13 <= _GEN_14;
                                                end else begin
                                                  if (6'hd == _T_218) begin
                                                    mem_13 <= _GEN_13;
                                                  end else begin
                                                    if (6'hd == _T_213) begin
                                                      mem_13 <= _GEN_12;
                                                    end else begin
                                                      if (6'hd == _T_208) begin
                                                        mem_13 <= _GEN_11;
                                                      end else begin
                                                        if (6'hd == _T_203) begin
                                                          mem_13 <= _GEN_10;
                                                        end else begin
                                                          if (6'hd == _T_198) begin
                                                            mem_13 <= _GEN_9;
                                                          end else begin
                                                            if (6'hd == _T_193) begin
                                                              mem_13 <= _GEN_8;
                                                            end else begin
                                                              if (6'hd == _T_188) begin
                                                                mem_13 <= _GEN_7;
                                                              end else begin
                                                                if (6'hd == _T_183) begin
                                                                  mem_13 <= _GEN_6;
                                                                end else begin
                                                                  if (6'hd == _T_178) begin
                                                                    mem_13 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'hd == _T_173) begin
                                                                      mem_13 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'hd == _T_168) begin
                                                                        mem_13 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'hd == _T_163) begin
                                                                          mem_13 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'hd == _T_158) begin
                                                                            mem_13 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'hd == _T_153) begin
                                                                              mem_13 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'hd == _T_308) begin
              mem_13 <= _GEN_31;
            end else begin
              if (6'hd == _T_303) begin
                mem_13 <= _GEN_30;
              end else begin
                if (6'hd == _T_298) begin
                  mem_13 <= _GEN_29;
                end else begin
                  if (6'hd == _T_293) begin
                    mem_13 <= _GEN_28;
                  end else begin
                    if (6'hd == _T_288) begin
                      mem_13 <= _GEN_27;
                    end else begin
                      if (6'hd == _T_283) begin
                        mem_13 <= _GEN_26;
                      end else begin
                        if (6'hd == _T_278) begin
                          mem_13 <= _GEN_25;
                        end else begin
                          if (6'hd == _T_273) begin
                            mem_13 <= _GEN_24;
                          end else begin
                            if (6'hd == _T_268) begin
                              mem_13 <= _GEN_23;
                            end else begin
                              if (6'hd == _T_263) begin
                                mem_13 <= _GEN_22;
                              end else begin
                                if (6'hd == _T_258) begin
                                  mem_13 <= _GEN_21;
                                end else begin
                                  if (6'hd == _T_253) begin
                                    mem_13 <= _GEN_20;
                                  end else begin
                                    if (6'hd == _T_248) begin
                                      mem_13 <= _GEN_19;
                                    end else begin
                                      if (6'hd == _T_243) begin
                                        mem_13 <= _GEN_18;
                                      end else begin
                                        if (6'hd == _T_238) begin
                                          mem_13 <= _GEN_17;
                                        end else begin
                                          if (6'hd == _T_233) begin
                                            mem_13 <= _GEN_16;
                                          end else begin
                                            if (6'hd == _T_228) begin
                                              mem_13 <= _GEN_15;
                                            end else begin
                                              if (6'hd == _T_223) begin
                                                mem_13 <= _GEN_14;
                                              end else begin
                                                if (6'hd == _T_218) begin
                                                  mem_13 <= _GEN_13;
                                                end else begin
                                                  if (6'hd == _T_213) begin
                                                    mem_13 <= _GEN_12;
                                                  end else begin
                                                    if (6'hd == _T_208) begin
                                                      mem_13 <= _GEN_11;
                                                    end else begin
                                                      if (6'hd == _T_203) begin
                                                        mem_13 <= _GEN_10;
                                                      end else begin
                                                        if (6'hd == _T_198) begin
                                                          mem_13 <= _GEN_9;
                                                        end else begin
                                                          if (6'hd == _T_193) begin
                                                            mem_13 <= _GEN_8;
                                                          end else begin
                                                            if (6'hd == _T_188) begin
                                                              mem_13 <= _GEN_7;
                                                            end else begin
                                                              if (6'hd == _T_183) begin
                                                                mem_13 <= _GEN_6;
                                                              end else begin
                                                                if (6'hd == _T_178) begin
                                                                  mem_13 <= _GEN_5;
                                                                end else begin
                                                                  if (6'hd == _T_173) begin
                                                                    mem_13 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'hd == _T_168) begin
                                                                      mem_13 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'hd == _T_163) begin
                                                                        mem_13 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'hd == _T_158) begin
                                                                          mem_13 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'hd == _T_153) begin
                                                                            mem_13 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'hd == _T_308) begin
            mem_13 <= _GEN_31;
          end else begin
            if (6'hd == _T_303) begin
              mem_13 <= _GEN_30;
            end else begin
              if (6'hd == _T_298) begin
                mem_13 <= _GEN_29;
              end else begin
                if (6'hd == _T_293) begin
                  mem_13 <= _GEN_28;
                end else begin
                  if (6'hd == _T_288) begin
                    mem_13 <= _GEN_27;
                  end else begin
                    if (6'hd == _T_283) begin
                      mem_13 <= _GEN_26;
                    end else begin
                      if (6'hd == _T_278) begin
                        mem_13 <= _GEN_25;
                      end else begin
                        if (6'hd == _T_273) begin
                          mem_13 <= _GEN_24;
                        end else begin
                          if (6'hd == _T_268) begin
                            mem_13 <= _GEN_23;
                          end else begin
                            if (6'hd == _T_263) begin
                              mem_13 <= _GEN_22;
                            end else begin
                              if (6'hd == _T_258) begin
                                mem_13 <= _GEN_21;
                              end else begin
                                if (6'hd == _T_253) begin
                                  mem_13 <= _GEN_20;
                                end else begin
                                  if (6'hd == _T_248) begin
                                    mem_13 <= _GEN_19;
                                  end else begin
                                    if (6'hd == _T_243) begin
                                      mem_13 <= _GEN_18;
                                    end else begin
                                      if (6'hd == _T_238) begin
                                        mem_13 <= _GEN_17;
                                      end else begin
                                        if (6'hd == _T_233) begin
                                          mem_13 <= _GEN_16;
                                        end else begin
                                          if (6'hd == _T_228) begin
                                            mem_13 <= _GEN_15;
                                          end else begin
                                            if (6'hd == _T_223) begin
                                              mem_13 <= _GEN_14;
                                            end else begin
                                              if (6'hd == _T_218) begin
                                                mem_13 <= _GEN_13;
                                              end else begin
                                                if (6'hd == _T_213) begin
                                                  mem_13 <= _GEN_12;
                                                end else begin
                                                  if (6'hd == _T_208) begin
                                                    mem_13 <= _GEN_11;
                                                  end else begin
                                                    if (6'hd == _T_203) begin
                                                      mem_13 <= _GEN_10;
                                                    end else begin
                                                      if (6'hd == _T_198) begin
                                                        mem_13 <= _GEN_9;
                                                      end else begin
                                                        if (6'hd == _T_193) begin
                                                          mem_13 <= _GEN_8;
                                                        end else begin
                                                          if (6'hd == _T_188) begin
                                                            mem_13 <= _GEN_7;
                                                          end else begin
                                                            if (6'hd == _T_183) begin
                                                              mem_13 <= _GEN_6;
                                                            end else begin
                                                              if (6'hd == _T_178) begin
                                                                mem_13 <= _GEN_5;
                                                              end else begin
                                                                if (6'hd == _T_173) begin
                                                                  mem_13 <= _GEN_4;
                                                                end else begin
                                                                  if (6'hd == _T_168) begin
                                                                    mem_13 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'hd == _T_163) begin
                                                                      mem_13 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'hd == _T_158) begin
                                                                        mem_13 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'hd == _T_153) begin
                                                                          mem_13 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'hd == _T_308) begin
          mem_13 <= _GEN_31;
        end else begin
          if (6'hd == _T_303) begin
            mem_13 <= _GEN_30;
          end else begin
            if (6'hd == _T_298) begin
              mem_13 <= _GEN_29;
            end else begin
              if (6'hd == _T_293) begin
                mem_13 <= _GEN_28;
              end else begin
                if (6'hd == _T_288) begin
                  mem_13 <= _GEN_27;
                end else begin
                  if (6'hd == _T_283) begin
                    mem_13 <= _GEN_26;
                  end else begin
                    if (6'hd == _T_278) begin
                      mem_13 <= _GEN_25;
                    end else begin
                      if (6'hd == _T_273) begin
                        mem_13 <= _GEN_24;
                      end else begin
                        if (6'hd == _T_268) begin
                          mem_13 <= _GEN_23;
                        end else begin
                          if (6'hd == _T_263) begin
                            mem_13 <= _GEN_22;
                          end else begin
                            if (6'hd == _T_258) begin
                              mem_13 <= _GEN_21;
                            end else begin
                              if (6'hd == _T_253) begin
                                mem_13 <= _GEN_20;
                              end else begin
                                if (6'hd == _T_248) begin
                                  mem_13 <= _GEN_19;
                                end else begin
                                  if (6'hd == _T_243) begin
                                    mem_13 <= _GEN_18;
                                  end else begin
                                    if (6'hd == _T_238) begin
                                      mem_13 <= _GEN_17;
                                    end else begin
                                      if (6'hd == _T_233) begin
                                        mem_13 <= _GEN_16;
                                      end else begin
                                        if (6'hd == _T_228) begin
                                          mem_13 <= _GEN_15;
                                        end else begin
                                          if (6'hd == _T_223) begin
                                            mem_13 <= _GEN_14;
                                          end else begin
                                            if (6'hd == _T_218) begin
                                              mem_13 <= _GEN_13;
                                            end else begin
                                              if (6'hd == _T_213) begin
                                                mem_13 <= _GEN_12;
                                              end else begin
                                                if (6'hd == _T_208) begin
                                                  mem_13 <= _GEN_11;
                                                end else begin
                                                  if (6'hd == _T_203) begin
                                                    mem_13 <= _GEN_10;
                                                  end else begin
                                                    if (6'hd == _T_198) begin
                                                      mem_13 <= _GEN_9;
                                                    end else begin
                                                      if (6'hd == _T_193) begin
                                                        mem_13 <= _GEN_8;
                                                      end else begin
                                                        if (6'hd == _T_188) begin
                                                          mem_13 <= _GEN_7;
                                                        end else begin
                                                          if (6'hd == _T_183) begin
                                                            mem_13 <= _GEN_6;
                                                          end else begin
                                                            if (6'hd == _T_178) begin
                                                              mem_13 <= _GEN_5;
                                                            end else begin
                                                              if (6'hd == _T_173) begin
                                                                mem_13 <= _GEN_4;
                                                              end else begin
                                                                if (6'hd == _T_168) begin
                                                                  mem_13 <= _GEN_3;
                                                                end else begin
                                                                  if (6'hd == _T_163) begin
                                                                    mem_13 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'hd == _T_158) begin
                                                                      mem_13 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'hd == _T_153) begin
                                                                        mem_13 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'he == wPos) begin
            mem_14 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'he == _T_308) begin
                mem_14 <= _GEN_31;
              end else begin
                if (6'he == _T_303) begin
                  mem_14 <= _GEN_30;
                end else begin
                  if (6'he == _T_298) begin
                    mem_14 <= _GEN_29;
                  end else begin
                    if (6'he == _T_293) begin
                      mem_14 <= _GEN_28;
                    end else begin
                      if (6'he == _T_288) begin
                        mem_14 <= _GEN_27;
                      end else begin
                        if (6'he == _T_283) begin
                          mem_14 <= _GEN_26;
                        end else begin
                          if (6'he == _T_278) begin
                            mem_14 <= _GEN_25;
                          end else begin
                            if (6'he == _T_273) begin
                              mem_14 <= _GEN_24;
                            end else begin
                              if (6'he == _T_268) begin
                                mem_14 <= _GEN_23;
                              end else begin
                                if (6'he == _T_263) begin
                                  mem_14 <= _GEN_22;
                                end else begin
                                  if (6'he == _T_258) begin
                                    mem_14 <= _GEN_21;
                                  end else begin
                                    if (6'he == _T_253) begin
                                      mem_14 <= _GEN_20;
                                    end else begin
                                      if (6'he == _T_248) begin
                                        mem_14 <= _GEN_19;
                                      end else begin
                                        if (6'he == _T_243) begin
                                          mem_14 <= _GEN_18;
                                        end else begin
                                          if (6'he == _T_238) begin
                                            mem_14 <= _GEN_17;
                                          end else begin
                                            if (6'he == _T_233) begin
                                              mem_14 <= _GEN_16;
                                            end else begin
                                              if (6'he == _T_228) begin
                                                mem_14 <= _GEN_15;
                                              end else begin
                                                if (6'he == _T_223) begin
                                                  mem_14 <= _GEN_14;
                                                end else begin
                                                  if (6'he == _T_218) begin
                                                    mem_14 <= _GEN_13;
                                                  end else begin
                                                    if (6'he == _T_213) begin
                                                      mem_14 <= _GEN_12;
                                                    end else begin
                                                      if (6'he == _T_208) begin
                                                        mem_14 <= _GEN_11;
                                                      end else begin
                                                        if (6'he == _T_203) begin
                                                          mem_14 <= _GEN_10;
                                                        end else begin
                                                          if (6'he == _T_198) begin
                                                            mem_14 <= _GEN_9;
                                                          end else begin
                                                            if (6'he == _T_193) begin
                                                              mem_14 <= _GEN_8;
                                                            end else begin
                                                              if (6'he == _T_188) begin
                                                                mem_14 <= _GEN_7;
                                                              end else begin
                                                                if (6'he == _T_183) begin
                                                                  mem_14 <= _GEN_6;
                                                                end else begin
                                                                  if (6'he == _T_178) begin
                                                                    mem_14 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'he == _T_173) begin
                                                                      mem_14 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'he == _T_168) begin
                                                                        mem_14 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'he == _T_163) begin
                                                                          mem_14 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'he == _T_158) begin
                                                                            mem_14 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'he == _T_153) begin
                                                                              mem_14 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'he == _T_308) begin
              mem_14 <= _GEN_31;
            end else begin
              if (6'he == _T_303) begin
                mem_14 <= _GEN_30;
              end else begin
                if (6'he == _T_298) begin
                  mem_14 <= _GEN_29;
                end else begin
                  if (6'he == _T_293) begin
                    mem_14 <= _GEN_28;
                  end else begin
                    if (6'he == _T_288) begin
                      mem_14 <= _GEN_27;
                    end else begin
                      if (6'he == _T_283) begin
                        mem_14 <= _GEN_26;
                      end else begin
                        if (6'he == _T_278) begin
                          mem_14 <= _GEN_25;
                        end else begin
                          if (6'he == _T_273) begin
                            mem_14 <= _GEN_24;
                          end else begin
                            if (6'he == _T_268) begin
                              mem_14 <= _GEN_23;
                            end else begin
                              if (6'he == _T_263) begin
                                mem_14 <= _GEN_22;
                              end else begin
                                if (6'he == _T_258) begin
                                  mem_14 <= _GEN_21;
                                end else begin
                                  if (6'he == _T_253) begin
                                    mem_14 <= _GEN_20;
                                  end else begin
                                    if (6'he == _T_248) begin
                                      mem_14 <= _GEN_19;
                                    end else begin
                                      if (6'he == _T_243) begin
                                        mem_14 <= _GEN_18;
                                      end else begin
                                        if (6'he == _T_238) begin
                                          mem_14 <= _GEN_17;
                                        end else begin
                                          if (6'he == _T_233) begin
                                            mem_14 <= _GEN_16;
                                          end else begin
                                            if (6'he == _T_228) begin
                                              mem_14 <= _GEN_15;
                                            end else begin
                                              if (6'he == _T_223) begin
                                                mem_14 <= _GEN_14;
                                              end else begin
                                                if (6'he == _T_218) begin
                                                  mem_14 <= _GEN_13;
                                                end else begin
                                                  if (6'he == _T_213) begin
                                                    mem_14 <= _GEN_12;
                                                  end else begin
                                                    if (6'he == _T_208) begin
                                                      mem_14 <= _GEN_11;
                                                    end else begin
                                                      if (6'he == _T_203) begin
                                                        mem_14 <= _GEN_10;
                                                      end else begin
                                                        if (6'he == _T_198) begin
                                                          mem_14 <= _GEN_9;
                                                        end else begin
                                                          if (6'he == _T_193) begin
                                                            mem_14 <= _GEN_8;
                                                          end else begin
                                                            if (6'he == _T_188) begin
                                                              mem_14 <= _GEN_7;
                                                            end else begin
                                                              if (6'he == _T_183) begin
                                                                mem_14 <= _GEN_6;
                                                              end else begin
                                                                if (6'he == _T_178) begin
                                                                  mem_14 <= _GEN_5;
                                                                end else begin
                                                                  if (6'he == _T_173) begin
                                                                    mem_14 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'he == _T_168) begin
                                                                      mem_14 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'he == _T_163) begin
                                                                        mem_14 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'he == _T_158) begin
                                                                          mem_14 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'he == _T_153) begin
                                                                            mem_14 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'he == _T_308) begin
            mem_14 <= _GEN_31;
          end else begin
            if (6'he == _T_303) begin
              mem_14 <= _GEN_30;
            end else begin
              if (6'he == _T_298) begin
                mem_14 <= _GEN_29;
              end else begin
                if (6'he == _T_293) begin
                  mem_14 <= _GEN_28;
                end else begin
                  if (6'he == _T_288) begin
                    mem_14 <= _GEN_27;
                  end else begin
                    if (6'he == _T_283) begin
                      mem_14 <= _GEN_26;
                    end else begin
                      if (6'he == _T_278) begin
                        mem_14 <= _GEN_25;
                      end else begin
                        if (6'he == _T_273) begin
                          mem_14 <= _GEN_24;
                        end else begin
                          if (6'he == _T_268) begin
                            mem_14 <= _GEN_23;
                          end else begin
                            if (6'he == _T_263) begin
                              mem_14 <= _GEN_22;
                            end else begin
                              if (6'he == _T_258) begin
                                mem_14 <= _GEN_21;
                              end else begin
                                if (6'he == _T_253) begin
                                  mem_14 <= _GEN_20;
                                end else begin
                                  if (6'he == _T_248) begin
                                    mem_14 <= _GEN_19;
                                  end else begin
                                    if (6'he == _T_243) begin
                                      mem_14 <= _GEN_18;
                                    end else begin
                                      if (6'he == _T_238) begin
                                        mem_14 <= _GEN_17;
                                      end else begin
                                        if (6'he == _T_233) begin
                                          mem_14 <= _GEN_16;
                                        end else begin
                                          if (6'he == _T_228) begin
                                            mem_14 <= _GEN_15;
                                          end else begin
                                            if (6'he == _T_223) begin
                                              mem_14 <= _GEN_14;
                                            end else begin
                                              if (6'he == _T_218) begin
                                                mem_14 <= _GEN_13;
                                              end else begin
                                                if (6'he == _T_213) begin
                                                  mem_14 <= _GEN_12;
                                                end else begin
                                                  if (6'he == _T_208) begin
                                                    mem_14 <= _GEN_11;
                                                  end else begin
                                                    if (6'he == _T_203) begin
                                                      mem_14 <= _GEN_10;
                                                    end else begin
                                                      if (6'he == _T_198) begin
                                                        mem_14 <= _GEN_9;
                                                      end else begin
                                                        if (6'he == _T_193) begin
                                                          mem_14 <= _GEN_8;
                                                        end else begin
                                                          if (6'he == _T_188) begin
                                                            mem_14 <= _GEN_7;
                                                          end else begin
                                                            if (6'he == _T_183) begin
                                                              mem_14 <= _GEN_6;
                                                            end else begin
                                                              if (6'he == _T_178) begin
                                                                mem_14 <= _GEN_5;
                                                              end else begin
                                                                if (6'he == _T_173) begin
                                                                  mem_14 <= _GEN_4;
                                                                end else begin
                                                                  if (6'he == _T_168) begin
                                                                    mem_14 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'he == _T_163) begin
                                                                      mem_14 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'he == _T_158) begin
                                                                        mem_14 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'he == _T_153) begin
                                                                          mem_14 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'he == _T_308) begin
          mem_14 <= _GEN_31;
        end else begin
          if (6'he == _T_303) begin
            mem_14 <= _GEN_30;
          end else begin
            if (6'he == _T_298) begin
              mem_14 <= _GEN_29;
            end else begin
              if (6'he == _T_293) begin
                mem_14 <= _GEN_28;
              end else begin
                if (6'he == _T_288) begin
                  mem_14 <= _GEN_27;
                end else begin
                  if (6'he == _T_283) begin
                    mem_14 <= _GEN_26;
                  end else begin
                    if (6'he == _T_278) begin
                      mem_14 <= _GEN_25;
                    end else begin
                      if (6'he == _T_273) begin
                        mem_14 <= _GEN_24;
                      end else begin
                        if (6'he == _T_268) begin
                          mem_14 <= _GEN_23;
                        end else begin
                          if (6'he == _T_263) begin
                            mem_14 <= _GEN_22;
                          end else begin
                            if (6'he == _T_258) begin
                              mem_14 <= _GEN_21;
                            end else begin
                              if (6'he == _T_253) begin
                                mem_14 <= _GEN_20;
                              end else begin
                                if (6'he == _T_248) begin
                                  mem_14 <= _GEN_19;
                                end else begin
                                  if (6'he == _T_243) begin
                                    mem_14 <= _GEN_18;
                                  end else begin
                                    if (6'he == _T_238) begin
                                      mem_14 <= _GEN_17;
                                    end else begin
                                      if (6'he == _T_233) begin
                                        mem_14 <= _GEN_16;
                                      end else begin
                                        if (6'he == _T_228) begin
                                          mem_14 <= _GEN_15;
                                        end else begin
                                          if (6'he == _T_223) begin
                                            mem_14 <= _GEN_14;
                                          end else begin
                                            if (6'he == _T_218) begin
                                              mem_14 <= _GEN_13;
                                            end else begin
                                              if (6'he == _T_213) begin
                                                mem_14 <= _GEN_12;
                                              end else begin
                                                if (6'he == _T_208) begin
                                                  mem_14 <= _GEN_11;
                                                end else begin
                                                  if (6'he == _T_203) begin
                                                    mem_14 <= _GEN_10;
                                                  end else begin
                                                    if (6'he == _T_198) begin
                                                      mem_14 <= _GEN_9;
                                                    end else begin
                                                      if (6'he == _T_193) begin
                                                        mem_14 <= _GEN_8;
                                                      end else begin
                                                        if (6'he == _T_188) begin
                                                          mem_14 <= _GEN_7;
                                                        end else begin
                                                          if (6'he == _T_183) begin
                                                            mem_14 <= _GEN_6;
                                                          end else begin
                                                            if (6'he == _T_178) begin
                                                              mem_14 <= _GEN_5;
                                                            end else begin
                                                              if (6'he == _T_173) begin
                                                                mem_14 <= _GEN_4;
                                                              end else begin
                                                                if (6'he == _T_168) begin
                                                                  mem_14 <= _GEN_3;
                                                                end else begin
                                                                  if (6'he == _T_163) begin
                                                                    mem_14 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'he == _T_158) begin
                                                                      mem_14 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'he == _T_153) begin
                                                                        mem_14 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'hf == wPos) begin
            mem_15 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'hf == _T_308) begin
                mem_15 <= _GEN_31;
              end else begin
                if (6'hf == _T_303) begin
                  mem_15 <= _GEN_30;
                end else begin
                  if (6'hf == _T_298) begin
                    mem_15 <= _GEN_29;
                  end else begin
                    if (6'hf == _T_293) begin
                      mem_15 <= _GEN_28;
                    end else begin
                      if (6'hf == _T_288) begin
                        mem_15 <= _GEN_27;
                      end else begin
                        if (6'hf == _T_283) begin
                          mem_15 <= _GEN_26;
                        end else begin
                          if (6'hf == _T_278) begin
                            mem_15 <= _GEN_25;
                          end else begin
                            if (6'hf == _T_273) begin
                              mem_15 <= _GEN_24;
                            end else begin
                              if (6'hf == _T_268) begin
                                mem_15 <= _GEN_23;
                              end else begin
                                if (6'hf == _T_263) begin
                                  mem_15 <= _GEN_22;
                                end else begin
                                  if (6'hf == _T_258) begin
                                    mem_15 <= _GEN_21;
                                  end else begin
                                    if (6'hf == _T_253) begin
                                      mem_15 <= _GEN_20;
                                    end else begin
                                      if (6'hf == _T_248) begin
                                        mem_15 <= _GEN_19;
                                      end else begin
                                        if (6'hf == _T_243) begin
                                          mem_15 <= _GEN_18;
                                        end else begin
                                          if (6'hf == _T_238) begin
                                            mem_15 <= _GEN_17;
                                          end else begin
                                            if (6'hf == _T_233) begin
                                              mem_15 <= _GEN_16;
                                            end else begin
                                              if (6'hf == _T_228) begin
                                                mem_15 <= _GEN_15;
                                              end else begin
                                                if (6'hf == _T_223) begin
                                                  mem_15 <= _GEN_14;
                                                end else begin
                                                  if (6'hf == _T_218) begin
                                                    mem_15 <= _GEN_13;
                                                  end else begin
                                                    if (6'hf == _T_213) begin
                                                      mem_15 <= _GEN_12;
                                                    end else begin
                                                      if (6'hf == _T_208) begin
                                                        mem_15 <= _GEN_11;
                                                      end else begin
                                                        if (6'hf == _T_203) begin
                                                          mem_15 <= _GEN_10;
                                                        end else begin
                                                          if (6'hf == _T_198) begin
                                                            mem_15 <= _GEN_9;
                                                          end else begin
                                                            if (6'hf == _T_193) begin
                                                              mem_15 <= _GEN_8;
                                                            end else begin
                                                              if (6'hf == _T_188) begin
                                                                mem_15 <= _GEN_7;
                                                              end else begin
                                                                if (6'hf == _T_183) begin
                                                                  mem_15 <= _GEN_6;
                                                                end else begin
                                                                  if (6'hf == _T_178) begin
                                                                    mem_15 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'hf == _T_173) begin
                                                                      mem_15 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'hf == _T_168) begin
                                                                        mem_15 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'hf == _T_163) begin
                                                                          mem_15 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'hf == _T_158) begin
                                                                            mem_15 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'hf == _T_153) begin
                                                                              mem_15 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'hf == _T_308) begin
              mem_15 <= _GEN_31;
            end else begin
              if (6'hf == _T_303) begin
                mem_15 <= _GEN_30;
              end else begin
                if (6'hf == _T_298) begin
                  mem_15 <= _GEN_29;
                end else begin
                  if (6'hf == _T_293) begin
                    mem_15 <= _GEN_28;
                  end else begin
                    if (6'hf == _T_288) begin
                      mem_15 <= _GEN_27;
                    end else begin
                      if (6'hf == _T_283) begin
                        mem_15 <= _GEN_26;
                      end else begin
                        if (6'hf == _T_278) begin
                          mem_15 <= _GEN_25;
                        end else begin
                          if (6'hf == _T_273) begin
                            mem_15 <= _GEN_24;
                          end else begin
                            if (6'hf == _T_268) begin
                              mem_15 <= _GEN_23;
                            end else begin
                              if (6'hf == _T_263) begin
                                mem_15 <= _GEN_22;
                              end else begin
                                if (6'hf == _T_258) begin
                                  mem_15 <= _GEN_21;
                                end else begin
                                  if (6'hf == _T_253) begin
                                    mem_15 <= _GEN_20;
                                  end else begin
                                    if (6'hf == _T_248) begin
                                      mem_15 <= _GEN_19;
                                    end else begin
                                      if (6'hf == _T_243) begin
                                        mem_15 <= _GEN_18;
                                      end else begin
                                        if (6'hf == _T_238) begin
                                          mem_15 <= _GEN_17;
                                        end else begin
                                          if (6'hf == _T_233) begin
                                            mem_15 <= _GEN_16;
                                          end else begin
                                            if (6'hf == _T_228) begin
                                              mem_15 <= _GEN_15;
                                            end else begin
                                              if (6'hf == _T_223) begin
                                                mem_15 <= _GEN_14;
                                              end else begin
                                                if (6'hf == _T_218) begin
                                                  mem_15 <= _GEN_13;
                                                end else begin
                                                  if (6'hf == _T_213) begin
                                                    mem_15 <= _GEN_12;
                                                  end else begin
                                                    if (6'hf == _T_208) begin
                                                      mem_15 <= _GEN_11;
                                                    end else begin
                                                      if (6'hf == _T_203) begin
                                                        mem_15 <= _GEN_10;
                                                      end else begin
                                                        if (6'hf == _T_198) begin
                                                          mem_15 <= _GEN_9;
                                                        end else begin
                                                          if (6'hf == _T_193) begin
                                                            mem_15 <= _GEN_8;
                                                          end else begin
                                                            if (6'hf == _T_188) begin
                                                              mem_15 <= _GEN_7;
                                                            end else begin
                                                              if (6'hf == _T_183) begin
                                                                mem_15 <= _GEN_6;
                                                              end else begin
                                                                if (6'hf == _T_178) begin
                                                                  mem_15 <= _GEN_5;
                                                                end else begin
                                                                  if (6'hf == _T_173) begin
                                                                    mem_15 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'hf == _T_168) begin
                                                                      mem_15 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'hf == _T_163) begin
                                                                        mem_15 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'hf == _T_158) begin
                                                                          mem_15 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'hf == _T_153) begin
                                                                            mem_15 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'hf == _T_308) begin
            mem_15 <= _GEN_31;
          end else begin
            if (6'hf == _T_303) begin
              mem_15 <= _GEN_30;
            end else begin
              if (6'hf == _T_298) begin
                mem_15 <= _GEN_29;
              end else begin
                if (6'hf == _T_293) begin
                  mem_15 <= _GEN_28;
                end else begin
                  if (6'hf == _T_288) begin
                    mem_15 <= _GEN_27;
                  end else begin
                    if (6'hf == _T_283) begin
                      mem_15 <= _GEN_26;
                    end else begin
                      if (6'hf == _T_278) begin
                        mem_15 <= _GEN_25;
                      end else begin
                        if (6'hf == _T_273) begin
                          mem_15 <= _GEN_24;
                        end else begin
                          if (6'hf == _T_268) begin
                            mem_15 <= _GEN_23;
                          end else begin
                            if (6'hf == _T_263) begin
                              mem_15 <= _GEN_22;
                            end else begin
                              if (6'hf == _T_258) begin
                                mem_15 <= _GEN_21;
                              end else begin
                                if (6'hf == _T_253) begin
                                  mem_15 <= _GEN_20;
                                end else begin
                                  if (6'hf == _T_248) begin
                                    mem_15 <= _GEN_19;
                                  end else begin
                                    if (6'hf == _T_243) begin
                                      mem_15 <= _GEN_18;
                                    end else begin
                                      if (6'hf == _T_238) begin
                                        mem_15 <= _GEN_17;
                                      end else begin
                                        if (6'hf == _T_233) begin
                                          mem_15 <= _GEN_16;
                                        end else begin
                                          if (6'hf == _T_228) begin
                                            mem_15 <= _GEN_15;
                                          end else begin
                                            if (6'hf == _T_223) begin
                                              mem_15 <= _GEN_14;
                                            end else begin
                                              if (6'hf == _T_218) begin
                                                mem_15 <= _GEN_13;
                                              end else begin
                                                if (6'hf == _T_213) begin
                                                  mem_15 <= _GEN_12;
                                                end else begin
                                                  if (6'hf == _T_208) begin
                                                    mem_15 <= _GEN_11;
                                                  end else begin
                                                    if (6'hf == _T_203) begin
                                                      mem_15 <= _GEN_10;
                                                    end else begin
                                                      if (6'hf == _T_198) begin
                                                        mem_15 <= _GEN_9;
                                                      end else begin
                                                        if (6'hf == _T_193) begin
                                                          mem_15 <= _GEN_8;
                                                        end else begin
                                                          if (6'hf == _T_188) begin
                                                            mem_15 <= _GEN_7;
                                                          end else begin
                                                            if (6'hf == _T_183) begin
                                                              mem_15 <= _GEN_6;
                                                            end else begin
                                                              if (6'hf == _T_178) begin
                                                                mem_15 <= _GEN_5;
                                                              end else begin
                                                                if (6'hf == _T_173) begin
                                                                  mem_15 <= _GEN_4;
                                                                end else begin
                                                                  if (6'hf == _T_168) begin
                                                                    mem_15 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'hf == _T_163) begin
                                                                      mem_15 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'hf == _T_158) begin
                                                                        mem_15 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'hf == _T_153) begin
                                                                          mem_15 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'hf == _T_308) begin
          mem_15 <= _GEN_31;
        end else begin
          if (6'hf == _T_303) begin
            mem_15 <= _GEN_30;
          end else begin
            if (6'hf == _T_298) begin
              mem_15 <= _GEN_29;
            end else begin
              if (6'hf == _T_293) begin
                mem_15 <= _GEN_28;
              end else begin
                if (6'hf == _T_288) begin
                  mem_15 <= _GEN_27;
                end else begin
                  if (6'hf == _T_283) begin
                    mem_15 <= _GEN_26;
                  end else begin
                    if (6'hf == _T_278) begin
                      mem_15 <= _GEN_25;
                    end else begin
                      if (6'hf == _T_273) begin
                        mem_15 <= _GEN_24;
                      end else begin
                        if (6'hf == _T_268) begin
                          mem_15 <= _GEN_23;
                        end else begin
                          if (6'hf == _T_263) begin
                            mem_15 <= _GEN_22;
                          end else begin
                            if (6'hf == _T_258) begin
                              mem_15 <= _GEN_21;
                            end else begin
                              if (6'hf == _T_253) begin
                                mem_15 <= _GEN_20;
                              end else begin
                                if (6'hf == _T_248) begin
                                  mem_15 <= _GEN_19;
                                end else begin
                                  if (6'hf == _T_243) begin
                                    mem_15 <= _GEN_18;
                                  end else begin
                                    if (6'hf == _T_238) begin
                                      mem_15 <= _GEN_17;
                                    end else begin
                                      if (6'hf == _T_233) begin
                                        mem_15 <= _GEN_16;
                                      end else begin
                                        if (6'hf == _T_228) begin
                                          mem_15 <= _GEN_15;
                                        end else begin
                                          if (6'hf == _T_223) begin
                                            mem_15 <= _GEN_14;
                                          end else begin
                                            if (6'hf == _T_218) begin
                                              mem_15 <= _GEN_13;
                                            end else begin
                                              if (6'hf == _T_213) begin
                                                mem_15 <= _GEN_12;
                                              end else begin
                                                if (6'hf == _T_208) begin
                                                  mem_15 <= _GEN_11;
                                                end else begin
                                                  if (6'hf == _T_203) begin
                                                    mem_15 <= _GEN_10;
                                                  end else begin
                                                    if (6'hf == _T_198) begin
                                                      mem_15 <= _GEN_9;
                                                    end else begin
                                                      if (6'hf == _T_193) begin
                                                        mem_15 <= _GEN_8;
                                                      end else begin
                                                        if (6'hf == _T_188) begin
                                                          mem_15 <= _GEN_7;
                                                        end else begin
                                                          if (6'hf == _T_183) begin
                                                            mem_15 <= _GEN_6;
                                                          end else begin
                                                            if (6'hf == _T_178) begin
                                                              mem_15 <= _GEN_5;
                                                            end else begin
                                                              if (6'hf == _T_173) begin
                                                                mem_15 <= _GEN_4;
                                                              end else begin
                                                                if (6'hf == _T_168) begin
                                                                  mem_15 <= _GEN_3;
                                                                end else begin
                                                                  if (6'hf == _T_163) begin
                                                                    mem_15 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'hf == _T_158) begin
                                                                      mem_15 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'hf == _T_153) begin
                                                                        mem_15 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h10 == wPos) begin
            mem_16 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h10 == _T_308) begin
                mem_16 <= _GEN_31;
              end else begin
                if (6'h10 == _T_303) begin
                  mem_16 <= _GEN_30;
                end else begin
                  if (6'h10 == _T_298) begin
                    mem_16 <= _GEN_29;
                  end else begin
                    if (6'h10 == _T_293) begin
                      mem_16 <= _GEN_28;
                    end else begin
                      if (6'h10 == _T_288) begin
                        mem_16 <= _GEN_27;
                      end else begin
                        if (6'h10 == _T_283) begin
                          mem_16 <= _GEN_26;
                        end else begin
                          if (6'h10 == _T_278) begin
                            mem_16 <= _GEN_25;
                          end else begin
                            if (6'h10 == _T_273) begin
                              mem_16 <= _GEN_24;
                            end else begin
                              if (6'h10 == _T_268) begin
                                mem_16 <= _GEN_23;
                              end else begin
                                if (6'h10 == _T_263) begin
                                  mem_16 <= _GEN_22;
                                end else begin
                                  if (6'h10 == _T_258) begin
                                    mem_16 <= _GEN_21;
                                  end else begin
                                    if (6'h10 == _T_253) begin
                                      mem_16 <= _GEN_20;
                                    end else begin
                                      if (6'h10 == _T_248) begin
                                        mem_16 <= _GEN_19;
                                      end else begin
                                        if (6'h10 == _T_243) begin
                                          mem_16 <= _GEN_18;
                                        end else begin
                                          if (6'h10 == _T_238) begin
                                            mem_16 <= _GEN_17;
                                          end else begin
                                            if (6'h10 == _T_233) begin
                                              mem_16 <= _GEN_16;
                                            end else begin
                                              if (6'h10 == _T_228) begin
                                                mem_16 <= _GEN_15;
                                              end else begin
                                                if (6'h10 == _T_223) begin
                                                  mem_16 <= _GEN_14;
                                                end else begin
                                                  if (6'h10 == _T_218) begin
                                                    mem_16 <= _GEN_13;
                                                  end else begin
                                                    if (6'h10 == _T_213) begin
                                                      mem_16 <= _GEN_12;
                                                    end else begin
                                                      if (6'h10 == _T_208) begin
                                                        mem_16 <= _GEN_11;
                                                      end else begin
                                                        if (6'h10 == _T_203) begin
                                                          mem_16 <= _GEN_10;
                                                        end else begin
                                                          if (6'h10 == _T_198) begin
                                                            mem_16 <= _GEN_9;
                                                          end else begin
                                                            if (6'h10 == _T_193) begin
                                                              mem_16 <= _GEN_8;
                                                            end else begin
                                                              if (6'h10 == _T_188) begin
                                                                mem_16 <= _GEN_7;
                                                              end else begin
                                                                if (6'h10 == _T_183) begin
                                                                  mem_16 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h10 == _T_178) begin
                                                                    mem_16 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h10 == _T_173) begin
                                                                      mem_16 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h10 == _T_168) begin
                                                                        mem_16 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h10 == _T_163) begin
                                                                          mem_16 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h10 == _T_158) begin
                                                                            mem_16 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h10 == _T_153) begin
                                                                              mem_16 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h10 == _T_308) begin
              mem_16 <= _GEN_31;
            end else begin
              if (6'h10 == _T_303) begin
                mem_16 <= _GEN_30;
              end else begin
                if (6'h10 == _T_298) begin
                  mem_16 <= _GEN_29;
                end else begin
                  if (6'h10 == _T_293) begin
                    mem_16 <= _GEN_28;
                  end else begin
                    if (6'h10 == _T_288) begin
                      mem_16 <= _GEN_27;
                    end else begin
                      if (6'h10 == _T_283) begin
                        mem_16 <= _GEN_26;
                      end else begin
                        if (6'h10 == _T_278) begin
                          mem_16 <= _GEN_25;
                        end else begin
                          if (6'h10 == _T_273) begin
                            mem_16 <= _GEN_24;
                          end else begin
                            if (6'h10 == _T_268) begin
                              mem_16 <= _GEN_23;
                            end else begin
                              if (6'h10 == _T_263) begin
                                mem_16 <= _GEN_22;
                              end else begin
                                if (6'h10 == _T_258) begin
                                  mem_16 <= _GEN_21;
                                end else begin
                                  if (6'h10 == _T_253) begin
                                    mem_16 <= _GEN_20;
                                  end else begin
                                    if (6'h10 == _T_248) begin
                                      mem_16 <= _GEN_19;
                                    end else begin
                                      if (6'h10 == _T_243) begin
                                        mem_16 <= _GEN_18;
                                      end else begin
                                        if (6'h10 == _T_238) begin
                                          mem_16 <= _GEN_17;
                                        end else begin
                                          if (6'h10 == _T_233) begin
                                            mem_16 <= _GEN_16;
                                          end else begin
                                            if (6'h10 == _T_228) begin
                                              mem_16 <= _GEN_15;
                                            end else begin
                                              if (6'h10 == _T_223) begin
                                                mem_16 <= _GEN_14;
                                              end else begin
                                                if (6'h10 == _T_218) begin
                                                  mem_16 <= _GEN_13;
                                                end else begin
                                                  if (6'h10 == _T_213) begin
                                                    mem_16 <= _GEN_12;
                                                  end else begin
                                                    if (6'h10 == _T_208) begin
                                                      mem_16 <= _GEN_11;
                                                    end else begin
                                                      if (6'h10 == _T_203) begin
                                                        mem_16 <= _GEN_10;
                                                      end else begin
                                                        if (6'h10 == _T_198) begin
                                                          mem_16 <= _GEN_9;
                                                        end else begin
                                                          if (6'h10 == _T_193) begin
                                                            mem_16 <= _GEN_8;
                                                          end else begin
                                                            if (6'h10 == _T_188) begin
                                                              mem_16 <= _GEN_7;
                                                            end else begin
                                                              if (6'h10 == _T_183) begin
                                                                mem_16 <= _GEN_6;
                                                              end else begin
                                                                if (6'h10 == _T_178) begin
                                                                  mem_16 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h10 == _T_173) begin
                                                                    mem_16 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h10 == _T_168) begin
                                                                      mem_16 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h10 == _T_163) begin
                                                                        mem_16 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h10 == _T_158) begin
                                                                          mem_16 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h10 == _T_153) begin
                                                                            mem_16 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h10 == _T_308) begin
            mem_16 <= _GEN_31;
          end else begin
            if (6'h10 == _T_303) begin
              mem_16 <= _GEN_30;
            end else begin
              if (6'h10 == _T_298) begin
                mem_16 <= _GEN_29;
              end else begin
                if (6'h10 == _T_293) begin
                  mem_16 <= _GEN_28;
                end else begin
                  if (6'h10 == _T_288) begin
                    mem_16 <= _GEN_27;
                  end else begin
                    if (6'h10 == _T_283) begin
                      mem_16 <= _GEN_26;
                    end else begin
                      if (6'h10 == _T_278) begin
                        mem_16 <= _GEN_25;
                      end else begin
                        if (6'h10 == _T_273) begin
                          mem_16 <= _GEN_24;
                        end else begin
                          if (6'h10 == _T_268) begin
                            mem_16 <= _GEN_23;
                          end else begin
                            if (6'h10 == _T_263) begin
                              mem_16 <= _GEN_22;
                            end else begin
                              if (6'h10 == _T_258) begin
                                mem_16 <= _GEN_21;
                              end else begin
                                if (6'h10 == _T_253) begin
                                  mem_16 <= _GEN_20;
                                end else begin
                                  if (6'h10 == _T_248) begin
                                    mem_16 <= _GEN_19;
                                  end else begin
                                    if (6'h10 == _T_243) begin
                                      mem_16 <= _GEN_18;
                                    end else begin
                                      if (6'h10 == _T_238) begin
                                        mem_16 <= _GEN_17;
                                      end else begin
                                        if (6'h10 == _T_233) begin
                                          mem_16 <= _GEN_16;
                                        end else begin
                                          if (6'h10 == _T_228) begin
                                            mem_16 <= _GEN_15;
                                          end else begin
                                            if (6'h10 == _T_223) begin
                                              mem_16 <= _GEN_14;
                                            end else begin
                                              if (6'h10 == _T_218) begin
                                                mem_16 <= _GEN_13;
                                              end else begin
                                                if (6'h10 == _T_213) begin
                                                  mem_16 <= _GEN_12;
                                                end else begin
                                                  if (6'h10 == _T_208) begin
                                                    mem_16 <= _GEN_11;
                                                  end else begin
                                                    if (6'h10 == _T_203) begin
                                                      mem_16 <= _GEN_10;
                                                    end else begin
                                                      if (6'h10 == _T_198) begin
                                                        mem_16 <= _GEN_9;
                                                      end else begin
                                                        if (6'h10 == _T_193) begin
                                                          mem_16 <= _GEN_8;
                                                        end else begin
                                                          if (6'h10 == _T_188) begin
                                                            mem_16 <= _GEN_7;
                                                          end else begin
                                                            if (6'h10 == _T_183) begin
                                                              mem_16 <= _GEN_6;
                                                            end else begin
                                                              if (6'h10 == _T_178) begin
                                                                mem_16 <= _GEN_5;
                                                              end else begin
                                                                if (6'h10 == _T_173) begin
                                                                  mem_16 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h10 == _T_168) begin
                                                                    mem_16 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h10 == _T_163) begin
                                                                      mem_16 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h10 == _T_158) begin
                                                                        mem_16 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h10 == _T_153) begin
                                                                          mem_16 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h10 == _T_308) begin
          mem_16 <= _GEN_31;
        end else begin
          if (6'h10 == _T_303) begin
            mem_16 <= _GEN_30;
          end else begin
            if (6'h10 == _T_298) begin
              mem_16 <= _GEN_29;
            end else begin
              if (6'h10 == _T_293) begin
                mem_16 <= _GEN_28;
              end else begin
                if (6'h10 == _T_288) begin
                  mem_16 <= _GEN_27;
                end else begin
                  if (6'h10 == _T_283) begin
                    mem_16 <= _GEN_26;
                  end else begin
                    if (6'h10 == _T_278) begin
                      mem_16 <= _GEN_25;
                    end else begin
                      if (6'h10 == _T_273) begin
                        mem_16 <= _GEN_24;
                      end else begin
                        if (6'h10 == _T_268) begin
                          mem_16 <= _GEN_23;
                        end else begin
                          if (6'h10 == _T_263) begin
                            mem_16 <= _GEN_22;
                          end else begin
                            if (6'h10 == _T_258) begin
                              mem_16 <= _GEN_21;
                            end else begin
                              if (6'h10 == _T_253) begin
                                mem_16 <= _GEN_20;
                              end else begin
                                if (6'h10 == _T_248) begin
                                  mem_16 <= _GEN_19;
                                end else begin
                                  if (6'h10 == _T_243) begin
                                    mem_16 <= _GEN_18;
                                  end else begin
                                    if (6'h10 == _T_238) begin
                                      mem_16 <= _GEN_17;
                                    end else begin
                                      if (6'h10 == _T_233) begin
                                        mem_16 <= _GEN_16;
                                      end else begin
                                        if (6'h10 == _T_228) begin
                                          mem_16 <= _GEN_15;
                                        end else begin
                                          if (6'h10 == _T_223) begin
                                            mem_16 <= _GEN_14;
                                          end else begin
                                            if (6'h10 == _T_218) begin
                                              mem_16 <= _GEN_13;
                                            end else begin
                                              if (6'h10 == _T_213) begin
                                                mem_16 <= _GEN_12;
                                              end else begin
                                                if (6'h10 == _T_208) begin
                                                  mem_16 <= _GEN_11;
                                                end else begin
                                                  if (6'h10 == _T_203) begin
                                                    mem_16 <= _GEN_10;
                                                  end else begin
                                                    if (6'h10 == _T_198) begin
                                                      mem_16 <= _GEN_9;
                                                    end else begin
                                                      if (6'h10 == _T_193) begin
                                                        mem_16 <= _GEN_8;
                                                      end else begin
                                                        if (6'h10 == _T_188) begin
                                                          mem_16 <= _GEN_7;
                                                        end else begin
                                                          if (6'h10 == _T_183) begin
                                                            mem_16 <= _GEN_6;
                                                          end else begin
                                                            if (6'h10 == _T_178) begin
                                                              mem_16 <= _GEN_5;
                                                            end else begin
                                                              if (6'h10 == _T_173) begin
                                                                mem_16 <= _GEN_4;
                                                              end else begin
                                                                if (6'h10 == _T_168) begin
                                                                  mem_16 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h10 == _T_163) begin
                                                                    mem_16 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h10 == _T_158) begin
                                                                      mem_16 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h10 == _T_153) begin
                                                                        mem_16 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h11 == wPos) begin
            mem_17 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h11 == _T_308) begin
                mem_17 <= _GEN_31;
              end else begin
                if (6'h11 == _T_303) begin
                  mem_17 <= _GEN_30;
                end else begin
                  if (6'h11 == _T_298) begin
                    mem_17 <= _GEN_29;
                  end else begin
                    if (6'h11 == _T_293) begin
                      mem_17 <= _GEN_28;
                    end else begin
                      if (6'h11 == _T_288) begin
                        mem_17 <= _GEN_27;
                      end else begin
                        if (6'h11 == _T_283) begin
                          mem_17 <= _GEN_26;
                        end else begin
                          if (6'h11 == _T_278) begin
                            mem_17 <= _GEN_25;
                          end else begin
                            if (6'h11 == _T_273) begin
                              mem_17 <= _GEN_24;
                            end else begin
                              if (6'h11 == _T_268) begin
                                mem_17 <= _GEN_23;
                              end else begin
                                if (6'h11 == _T_263) begin
                                  mem_17 <= _GEN_22;
                                end else begin
                                  if (6'h11 == _T_258) begin
                                    mem_17 <= _GEN_21;
                                  end else begin
                                    if (6'h11 == _T_253) begin
                                      mem_17 <= _GEN_20;
                                    end else begin
                                      if (6'h11 == _T_248) begin
                                        mem_17 <= _GEN_19;
                                      end else begin
                                        if (6'h11 == _T_243) begin
                                          mem_17 <= _GEN_18;
                                        end else begin
                                          if (6'h11 == _T_238) begin
                                            mem_17 <= _GEN_17;
                                          end else begin
                                            if (6'h11 == _T_233) begin
                                              mem_17 <= _GEN_16;
                                            end else begin
                                              if (6'h11 == _T_228) begin
                                                mem_17 <= _GEN_15;
                                              end else begin
                                                if (6'h11 == _T_223) begin
                                                  mem_17 <= _GEN_14;
                                                end else begin
                                                  if (6'h11 == _T_218) begin
                                                    mem_17 <= _GEN_13;
                                                  end else begin
                                                    if (6'h11 == _T_213) begin
                                                      mem_17 <= _GEN_12;
                                                    end else begin
                                                      if (6'h11 == _T_208) begin
                                                        mem_17 <= _GEN_11;
                                                      end else begin
                                                        if (6'h11 == _T_203) begin
                                                          mem_17 <= _GEN_10;
                                                        end else begin
                                                          if (6'h11 == _T_198) begin
                                                            mem_17 <= _GEN_9;
                                                          end else begin
                                                            if (6'h11 == _T_193) begin
                                                              mem_17 <= _GEN_8;
                                                            end else begin
                                                              if (6'h11 == _T_188) begin
                                                                mem_17 <= _GEN_7;
                                                              end else begin
                                                                if (6'h11 == _T_183) begin
                                                                  mem_17 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h11 == _T_178) begin
                                                                    mem_17 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h11 == _T_173) begin
                                                                      mem_17 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h11 == _T_168) begin
                                                                        mem_17 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h11 == _T_163) begin
                                                                          mem_17 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h11 == _T_158) begin
                                                                            mem_17 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h11 == _T_153) begin
                                                                              mem_17 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h11 == _T_308) begin
              mem_17 <= _GEN_31;
            end else begin
              if (6'h11 == _T_303) begin
                mem_17 <= _GEN_30;
              end else begin
                if (6'h11 == _T_298) begin
                  mem_17 <= _GEN_29;
                end else begin
                  if (6'h11 == _T_293) begin
                    mem_17 <= _GEN_28;
                  end else begin
                    if (6'h11 == _T_288) begin
                      mem_17 <= _GEN_27;
                    end else begin
                      if (6'h11 == _T_283) begin
                        mem_17 <= _GEN_26;
                      end else begin
                        if (6'h11 == _T_278) begin
                          mem_17 <= _GEN_25;
                        end else begin
                          if (6'h11 == _T_273) begin
                            mem_17 <= _GEN_24;
                          end else begin
                            if (6'h11 == _T_268) begin
                              mem_17 <= _GEN_23;
                            end else begin
                              if (6'h11 == _T_263) begin
                                mem_17 <= _GEN_22;
                              end else begin
                                if (6'h11 == _T_258) begin
                                  mem_17 <= _GEN_21;
                                end else begin
                                  if (6'h11 == _T_253) begin
                                    mem_17 <= _GEN_20;
                                  end else begin
                                    if (6'h11 == _T_248) begin
                                      mem_17 <= _GEN_19;
                                    end else begin
                                      if (6'h11 == _T_243) begin
                                        mem_17 <= _GEN_18;
                                      end else begin
                                        if (6'h11 == _T_238) begin
                                          mem_17 <= _GEN_17;
                                        end else begin
                                          if (6'h11 == _T_233) begin
                                            mem_17 <= _GEN_16;
                                          end else begin
                                            if (6'h11 == _T_228) begin
                                              mem_17 <= _GEN_15;
                                            end else begin
                                              if (6'h11 == _T_223) begin
                                                mem_17 <= _GEN_14;
                                              end else begin
                                                if (6'h11 == _T_218) begin
                                                  mem_17 <= _GEN_13;
                                                end else begin
                                                  if (6'h11 == _T_213) begin
                                                    mem_17 <= _GEN_12;
                                                  end else begin
                                                    if (6'h11 == _T_208) begin
                                                      mem_17 <= _GEN_11;
                                                    end else begin
                                                      if (6'h11 == _T_203) begin
                                                        mem_17 <= _GEN_10;
                                                      end else begin
                                                        if (6'h11 == _T_198) begin
                                                          mem_17 <= _GEN_9;
                                                        end else begin
                                                          if (6'h11 == _T_193) begin
                                                            mem_17 <= _GEN_8;
                                                          end else begin
                                                            if (6'h11 == _T_188) begin
                                                              mem_17 <= _GEN_7;
                                                            end else begin
                                                              if (6'h11 == _T_183) begin
                                                                mem_17 <= _GEN_6;
                                                              end else begin
                                                                if (6'h11 == _T_178) begin
                                                                  mem_17 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h11 == _T_173) begin
                                                                    mem_17 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h11 == _T_168) begin
                                                                      mem_17 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h11 == _T_163) begin
                                                                        mem_17 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h11 == _T_158) begin
                                                                          mem_17 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h11 == _T_153) begin
                                                                            mem_17 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h11 == _T_308) begin
            mem_17 <= _GEN_31;
          end else begin
            if (6'h11 == _T_303) begin
              mem_17 <= _GEN_30;
            end else begin
              if (6'h11 == _T_298) begin
                mem_17 <= _GEN_29;
              end else begin
                if (6'h11 == _T_293) begin
                  mem_17 <= _GEN_28;
                end else begin
                  if (6'h11 == _T_288) begin
                    mem_17 <= _GEN_27;
                  end else begin
                    if (6'h11 == _T_283) begin
                      mem_17 <= _GEN_26;
                    end else begin
                      if (6'h11 == _T_278) begin
                        mem_17 <= _GEN_25;
                      end else begin
                        if (6'h11 == _T_273) begin
                          mem_17 <= _GEN_24;
                        end else begin
                          if (6'h11 == _T_268) begin
                            mem_17 <= _GEN_23;
                          end else begin
                            if (6'h11 == _T_263) begin
                              mem_17 <= _GEN_22;
                            end else begin
                              if (6'h11 == _T_258) begin
                                mem_17 <= _GEN_21;
                              end else begin
                                if (6'h11 == _T_253) begin
                                  mem_17 <= _GEN_20;
                                end else begin
                                  if (6'h11 == _T_248) begin
                                    mem_17 <= _GEN_19;
                                  end else begin
                                    if (6'h11 == _T_243) begin
                                      mem_17 <= _GEN_18;
                                    end else begin
                                      if (6'h11 == _T_238) begin
                                        mem_17 <= _GEN_17;
                                      end else begin
                                        if (6'h11 == _T_233) begin
                                          mem_17 <= _GEN_16;
                                        end else begin
                                          if (6'h11 == _T_228) begin
                                            mem_17 <= _GEN_15;
                                          end else begin
                                            if (6'h11 == _T_223) begin
                                              mem_17 <= _GEN_14;
                                            end else begin
                                              if (6'h11 == _T_218) begin
                                                mem_17 <= _GEN_13;
                                              end else begin
                                                if (6'h11 == _T_213) begin
                                                  mem_17 <= _GEN_12;
                                                end else begin
                                                  if (6'h11 == _T_208) begin
                                                    mem_17 <= _GEN_11;
                                                  end else begin
                                                    if (6'h11 == _T_203) begin
                                                      mem_17 <= _GEN_10;
                                                    end else begin
                                                      if (6'h11 == _T_198) begin
                                                        mem_17 <= _GEN_9;
                                                      end else begin
                                                        if (6'h11 == _T_193) begin
                                                          mem_17 <= _GEN_8;
                                                        end else begin
                                                          if (6'h11 == _T_188) begin
                                                            mem_17 <= _GEN_7;
                                                          end else begin
                                                            if (6'h11 == _T_183) begin
                                                              mem_17 <= _GEN_6;
                                                            end else begin
                                                              if (6'h11 == _T_178) begin
                                                                mem_17 <= _GEN_5;
                                                              end else begin
                                                                if (6'h11 == _T_173) begin
                                                                  mem_17 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h11 == _T_168) begin
                                                                    mem_17 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h11 == _T_163) begin
                                                                      mem_17 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h11 == _T_158) begin
                                                                        mem_17 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h11 == _T_153) begin
                                                                          mem_17 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h11 == _T_308) begin
          mem_17 <= _GEN_31;
        end else begin
          if (6'h11 == _T_303) begin
            mem_17 <= _GEN_30;
          end else begin
            if (6'h11 == _T_298) begin
              mem_17 <= _GEN_29;
            end else begin
              if (6'h11 == _T_293) begin
                mem_17 <= _GEN_28;
              end else begin
                if (6'h11 == _T_288) begin
                  mem_17 <= _GEN_27;
                end else begin
                  if (6'h11 == _T_283) begin
                    mem_17 <= _GEN_26;
                  end else begin
                    if (6'h11 == _T_278) begin
                      mem_17 <= _GEN_25;
                    end else begin
                      if (6'h11 == _T_273) begin
                        mem_17 <= _GEN_24;
                      end else begin
                        if (6'h11 == _T_268) begin
                          mem_17 <= _GEN_23;
                        end else begin
                          if (6'h11 == _T_263) begin
                            mem_17 <= _GEN_22;
                          end else begin
                            if (6'h11 == _T_258) begin
                              mem_17 <= _GEN_21;
                            end else begin
                              if (6'h11 == _T_253) begin
                                mem_17 <= _GEN_20;
                              end else begin
                                if (6'h11 == _T_248) begin
                                  mem_17 <= _GEN_19;
                                end else begin
                                  if (6'h11 == _T_243) begin
                                    mem_17 <= _GEN_18;
                                  end else begin
                                    if (6'h11 == _T_238) begin
                                      mem_17 <= _GEN_17;
                                    end else begin
                                      if (6'h11 == _T_233) begin
                                        mem_17 <= _GEN_16;
                                      end else begin
                                        if (6'h11 == _T_228) begin
                                          mem_17 <= _GEN_15;
                                        end else begin
                                          if (6'h11 == _T_223) begin
                                            mem_17 <= _GEN_14;
                                          end else begin
                                            if (6'h11 == _T_218) begin
                                              mem_17 <= _GEN_13;
                                            end else begin
                                              if (6'h11 == _T_213) begin
                                                mem_17 <= _GEN_12;
                                              end else begin
                                                if (6'h11 == _T_208) begin
                                                  mem_17 <= _GEN_11;
                                                end else begin
                                                  if (6'h11 == _T_203) begin
                                                    mem_17 <= _GEN_10;
                                                  end else begin
                                                    if (6'h11 == _T_198) begin
                                                      mem_17 <= _GEN_9;
                                                    end else begin
                                                      if (6'h11 == _T_193) begin
                                                        mem_17 <= _GEN_8;
                                                      end else begin
                                                        if (6'h11 == _T_188) begin
                                                          mem_17 <= _GEN_7;
                                                        end else begin
                                                          if (6'h11 == _T_183) begin
                                                            mem_17 <= _GEN_6;
                                                          end else begin
                                                            if (6'h11 == _T_178) begin
                                                              mem_17 <= _GEN_5;
                                                            end else begin
                                                              if (6'h11 == _T_173) begin
                                                                mem_17 <= _GEN_4;
                                                              end else begin
                                                                if (6'h11 == _T_168) begin
                                                                  mem_17 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h11 == _T_163) begin
                                                                    mem_17 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h11 == _T_158) begin
                                                                      mem_17 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h11 == _T_153) begin
                                                                        mem_17 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h12 == wPos) begin
            mem_18 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h12 == _T_308) begin
                mem_18 <= _GEN_31;
              end else begin
                if (6'h12 == _T_303) begin
                  mem_18 <= _GEN_30;
                end else begin
                  if (6'h12 == _T_298) begin
                    mem_18 <= _GEN_29;
                  end else begin
                    if (6'h12 == _T_293) begin
                      mem_18 <= _GEN_28;
                    end else begin
                      if (6'h12 == _T_288) begin
                        mem_18 <= _GEN_27;
                      end else begin
                        if (6'h12 == _T_283) begin
                          mem_18 <= _GEN_26;
                        end else begin
                          if (6'h12 == _T_278) begin
                            mem_18 <= _GEN_25;
                          end else begin
                            if (6'h12 == _T_273) begin
                              mem_18 <= _GEN_24;
                            end else begin
                              if (6'h12 == _T_268) begin
                                mem_18 <= _GEN_23;
                              end else begin
                                if (6'h12 == _T_263) begin
                                  mem_18 <= _GEN_22;
                                end else begin
                                  if (6'h12 == _T_258) begin
                                    mem_18 <= _GEN_21;
                                  end else begin
                                    if (6'h12 == _T_253) begin
                                      mem_18 <= _GEN_20;
                                    end else begin
                                      if (6'h12 == _T_248) begin
                                        mem_18 <= _GEN_19;
                                      end else begin
                                        if (6'h12 == _T_243) begin
                                          mem_18 <= _GEN_18;
                                        end else begin
                                          if (6'h12 == _T_238) begin
                                            mem_18 <= _GEN_17;
                                          end else begin
                                            if (6'h12 == _T_233) begin
                                              mem_18 <= _GEN_16;
                                            end else begin
                                              if (6'h12 == _T_228) begin
                                                mem_18 <= _GEN_15;
                                              end else begin
                                                if (6'h12 == _T_223) begin
                                                  mem_18 <= _GEN_14;
                                                end else begin
                                                  if (6'h12 == _T_218) begin
                                                    mem_18 <= _GEN_13;
                                                  end else begin
                                                    if (6'h12 == _T_213) begin
                                                      mem_18 <= _GEN_12;
                                                    end else begin
                                                      if (6'h12 == _T_208) begin
                                                        mem_18 <= _GEN_11;
                                                      end else begin
                                                        if (6'h12 == _T_203) begin
                                                          mem_18 <= _GEN_10;
                                                        end else begin
                                                          if (6'h12 == _T_198) begin
                                                            mem_18 <= _GEN_9;
                                                          end else begin
                                                            if (6'h12 == _T_193) begin
                                                              mem_18 <= _GEN_8;
                                                            end else begin
                                                              if (6'h12 == _T_188) begin
                                                                mem_18 <= _GEN_7;
                                                              end else begin
                                                                if (6'h12 == _T_183) begin
                                                                  mem_18 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h12 == _T_178) begin
                                                                    mem_18 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h12 == _T_173) begin
                                                                      mem_18 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h12 == _T_168) begin
                                                                        mem_18 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h12 == _T_163) begin
                                                                          mem_18 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h12 == _T_158) begin
                                                                            mem_18 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h12 == _T_153) begin
                                                                              mem_18 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h12 == _T_308) begin
              mem_18 <= _GEN_31;
            end else begin
              if (6'h12 == _T_303) begin
                mem_18 <= _GEN_30;
              end else begin
                if (6'h12 == _T_298) begin
                  mem_18 <= _GEN_29;
                end else begin
                  if (6'h12 == _T_293) begin
                    mem_18 <= _GEN_28;
                  end else begin
                    if (6'h12 == _T_288) begin
                      mem_18 <= _GEN_27;
                    end else begin
                      if (6'h12 == _T_283) begin
                        mem_18 <= _GEN_26;
                      end else begin
                        if (6'h12 == _T_278) begin
                          mem_18 <= _GEN_25;
                        end else begin
                          if (6'h12 == _T_273) begin
                            mem_18 <= _GEN_24;
                          end else begin
                            if (6'h12 == _T_268) begin
                              mem_18 <= _GEN_23;
                            end else begin
                              if (6'h12 == _T_263) begin
                                mem_18 <= _GEN_22;
                              end else begin
                                if (6'h12 == _T_258) begin
                                  mem_18 <= _GEN_21;
                                end else begin
                                  if (6'h12 == _T_253) begin
                                    mem_18 <= _GEN_20;
                                  end else begin
                                    if (6'h12 == _T_248) begin
                                      mem_18 <= _GEN_19;
                                    end else begin
                                      if (6'h12 == _T_243) begin
                                        mem_18 <= _GEN_18;
                                      end else begin
                                        if (6'h12 == _T_238) begin
                                          mem_18 <= _GEN_17;
                                        end else begin
                                          if (6'h12 == _T_233) begin
                                            mem_18 <= _GEN_16;
                                          end else begin
                                            if (6'h12 == _T_228) begin
                                              mem_18 <= _GEN_15;
                                            end else begin
                                              if (6'h12 == _T_223) begin
                                                mem_18 <= _GEN_14;
                                              end else begin
                                                if (6'h12 == _T_218) begin
                                                  mem_18 <= _GEN_13;
                                                end else begin
                                                  if (6'h12 == _T_213) begin
                                                    mem_18 <= _GEN_12;
                                                  end else begin
                                                    if (6'h12 == _T_208) begin
                                                      mem_18 <= _GEN_11;
                                                    end else begin
                                                      if (6'h12 == _T_203) begin
                                                        mem_18 <= _GEN_10;
                                                      end else begin
                                                        if (6'h12 == _T_198) begin
                                                          mem_18 <= _GEN_9;
                                                        end else begin
                                                          if (6'h12 == _T_193) begin
                                                            mem_18 <= _GEN_8;
                                                          end else begin
                                                            if (6'h12 == _T_188) begin
                                                              mem_18 <= _GEN_7;
                                                            end else begin
                                                              if (6'h12 == _T_183) begin
                                                                mem_18 <= _GEN_6;
                                                              end else begin
                                                                if (6'h12 == _T_178) begin
                                                                  mem_18 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h12 == _T_173) begin
                                                                    mem_18 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h12 == _T_168) begin
                                                                      mem_18 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h12 == _T_163) begin
                                                                        mem_18 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h12 == _T_158) begin
                                                                          mem_18 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h12 == _T_153) begin
                                                                            mem_18 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h12 == _T_308) begin
            mem_18 <= _GEN_31;
          end else begin
            if (6'h12 == _T_303) begin
              mem_18 <= _GEN_30;
            end else begin
              if (6'h12 == _T_298) begin
                mem_18 <= _GEN_29;
              end else begin
                if (6'h12 == _T_293) begin
                  mem_18 <= _GEN_28;
                end else begin
                  if (6'h12 == _T_288) begin
                    mem_18 <= _GEN_27;
                  end else begin
                    if (6'h12 == _T_283) begin
                      mem_18 <= _GEN_26;
                    end else begin
                      if (6'h12 == _T_278) begin
                        mem_18 <= _GEN_25;
                      end else begin
                        if (6'h12 == _T_273) begin
                          mem_18 <= _GEN_24;
                        end else begin
                          if (6'h12 == _T_268) begin
                            mem_18 <= _GEN_23;
                          end else begin
                            if (6'h12 == _T_263) begin
                              mem_18 <= _GEN_22;
                            end else begin
                              if (6'h12 == _T_258) begin
                                mem_18 <= _GEN_21;
                              end else begin
                                if (6'h12 == _T_253) begin
                                  mem_18 <= _GEN_20;
                                end else begin
                                  if (6'h12 == _T_248) begin
                                    mem_18 <= _GEN_19;
                                  end else begin
                                    if (6'h12 == _T_243) begin
                                      mem_18 <= _GEN_18;
                                    end else begin
                                      if (6'h12 == _T_238) begin
                                        mem_18 <= _GEN_17;
                                      end else begin
                                        if (6'h12 == _T_233) begin
                                          mem_18 <= _GEN_16;
                                        end else begin
                                          if (6'h12 == _T_228) begin
                                            mem_18 <= _GEN_15;
                                          end else begin
                                            if (6'h12 == _T_223) begin
                                              mem_18 <= _GEN_14;
                                            end else begin
                                              if (6'h12 == _T_218) begin
                                                mem_18 <= _GEN_13;
                                              end else begin
                                                if (6'h12 == _T_213) begin
                                                  mem_18 <= _GEN_12;
                                                end else begin
                                                  if (6'h12 == _T_208) begin
                                                    mem_18 <= _GEN_11;
                                                  end else begin
                                                    if (6'h12 == _T_203) begin
                                                      mem_18 <= _GEN_10;
                                                    end else begin
                                                      if (6'h12 == _T_198) begin
                                                        mem_18 <= _GEN_9;
                                                      end else begin
                                                        if (6'h12 == _T_193) begin
                                                          mem_18 <= _GEN_8;
                                                        end else begin
                                                          if (6'h12 == _T_188) begin
                                                            mem_18 <= _GEN_7;
                                                          end else begin
                                                            if (6'h12 == _T_183) begin
                                                              mem_18 <= _GEN_6;
                                                            end else begin
                                                              if (6'h12 == _T_178) begin
                                                                mem_18 <= _GEN_5;
                                                              end else begin
                                                                if (6'h12 == _T_173) begin
                                                                  mem_18 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h12 == _T_168) begin
                                                                    mem_18 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h12 == _T_163) begin
                                                                      mem_18 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h12 == _T_158) begin
                                                                        mem_18 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h12 == _T_153) begin
                                                                          mem_18 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h12 == _T_308) begin
          mem_18 <= _GEN_31;
        end else begin
          if (6'h12 == _T_303) begin
            mem_18 <= _GEN_30;
          end else begin
            if (6'h12 == _T_298) begin
              mem_18 <= _GEN_29;
            end else begin
              if (6'h12 == _T_293) begin
                mem_18 <= _GEN_28;
              end else begin
                if (6'h12 == _T_288) begin
                  mem_18 <= _GEN_27;
                end else begin
                  if (6'h12 == _T_283) begin
                    mem_18 <= _GEN_26;
                  end else begin
                    if (6'h12 == _T_278) begin
                      mem_18 <= _GEN_25;
                    end else begin
                      if (6'h12 == _T_273) begin
                        mem_18 <= _GEN_24;
                      end else begin
                        if (6'h12 == _T_268) begin
                          mem_18 <= _GEN_23;
                        end else begin
                          if (6'h12 == _T_263) begin
                            mem_18 <= _GEN_22;
                          end else begin
                            if (6'h12 == _T_258) begin
                              mem_18 <= _GEN_21;
                            end else begin
                              if (6'h12 == _T_253) begin
                                mem_18 <= _GEN_20;
                              end else begin
                                if (6'h12 == _T_248) begin
                                  mem_18 <= _GEN_19;
                                end else begin
                                  if (6'h12 == _T_243) begin
                                    mem_18 <= _GEN_18;
                                  end else begin
                                    if (6'h12 == _T_238) begin
                                      mem_18 <= _GEN_17;
                                    end else begin
                                      if (6'h12 == _T_233) begin
                                        mem_18 <= _GEN_16;
                                      end else begin
                                        if (6'h12 == _T_228) begin
                                          mem_18 <= _GEN_15;
                                        end else begin
                                          if (6'h12 == _T_223) begin
                                            mem_18 <= _GEN_14;
                                          end else begin
                                            if (6'h12 == _T_218) begin
                                              mem_18 <= _GEN_13;
                                            end else begin
                                              if (6'h12 == _T_213) begin
                                                mem_18 <= _GEN_12;
                                              end else begin
                                                if (6'h12 == _T_208) begin
                                                  mem_18 <= _GEN_11;
                                                end else begin
                                                  if (6'h12 == _T_203) begin
                                                    mem_18 <= _GEN_10;
                                                  end else begin
                                                    if (6'h12 == _T_198) begin
                                                      mem_18 <= _GEN_9;
                                                    end else begin
                                                      if (6'h12 == _T_193) begin
                                                        mem_18 <= _GEN_8;
                                                      end else begin
                                                        if (6'h12 == _T_188) begin
                                                          mem_18 <= _GEN_7;
                                                        end else begin
                                                          if (6'h12 == _T_183) begin
                                                            mem_18 <= _GEN_6;
                                                          end else begin
                                                            if (6'h12 == _T_178) begin
                                                              mem_18 <= _GEN_5;
                                                            end else begin
                                                              if (6'h12 == _T_173) begin
                                                                mem_18 <= _GEN_4;
                                                              end else begin
                                                                if (6'h12 == _T_168) begin
                                                                  mem_18 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h12 == _T_163) begin
                                                                    mem_18 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h12 == _T_158) begin
                                                                      mem_18 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h12 == _T_153) begin
                                                                        mem_18 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h13 == wPos) begin
            mem_19 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h13 == _T_308) begin
                mem_19 <= _GEN_31;
              end else begin
                if (6'h13 == _T_303) begin
                  mem_19 <= _GEN_30;
                end else begin
                  if (6'h13 == _T_298) begin
                    mem_19 <= _GEN_29;
                  end else begin
                    if (6'h13 == _T_293) begin
                      mem_19 <= _GEN_28;
                    end else begin
                      if (6'h13 == _T_288) begin
                        mem_19 <= _GEN_27;
                      end else begin
                        if (6'h13 == _T_283) begin
                          mem_19 <= _GEN_26;
                        end else begin
                          if (6'h13 == _T_278) begin
                            mem_19 <= _GEN_25;
                          end else begin
                            if (6'h13 == _T_273) begin
                              mem_19 <= _GEN_24;
                            end else begin
                              if (6'h13 == _T_268) begin
                                mem_19 <= _GEN_23;
                              end else begin
                                if (6'h13 == _T_263) begin
                                  mem_19 <= _GEN_22;
                                end else begin
                                  if (6'h13 == _T_258) begin
                                    mem_19 <= _GEN_21;
                                  end else begin
                                    if (6'h13 == _T_253) begin
                                      mem_19 <= _GEN_20;
                                    end else begin
                                      if (6'h13 == _T_248) begin
                                        mem_19 <= _GEN_19;
                                      end else begin
                                        if (6'h13 == _T_243) begin
                                          mem_19 <= _GEN_18;
                                        end else begin
                                          if (6'h13 == _T_238) begin
                                            mem_19 <= _GEN_17;
                                          end else begin
                                            if (6'h13 == _T_233) begin
                                              mem_19 <= _GEN_16;
                                            end else begin
                                              if (6'h13 == _T_228) begin
                                                mem_19 <= _GEN_15;
                                              end else begin
                                                if (6'h13 == _T_223) begin
                                                  mem_19 <= _GEN_14;
                                                end else begin
                                                  if (6'h13 == _T_218) begin
                                                    mem_19 <= _GEN_13;
                                                  end else begin
                                                    if (6'h13 == _T_213) begin
                                                      mem_19 <= _GEN_12;
                                                    end else begin
                                                      if (6'h13 == _T_208) begin
                                                        mem_19 <= _GEN_11;
                                                      end else begin
                                                        if (6'h13 == _T_203) begin
                                                          mem_19 <= _GEN_10;
                                                        end else begin
                                                          if (6'h13 == _T_198) begin
                                                            mem_19 <= _GEN_9;
                                                          end else begin
                                                            if (6'h13 == _T_193) begin
                                                              mem_19 <= _GEN_8;
                                                            end else begin
                                                              if (6'h13 == _T_188) begin
                                                                mem_19 <= _GEN_7;
                                                              end else begin
                                                                if (6'h13 == _T_183) begin
                                                                  mem_19 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h13 == _T_178) begin
                                                                    mem_19 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h13 == _T_173) begin
                                                                      mem_19 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h13 == _T_168) begin
                                                                        mem_19 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h13 == _T_163) begin
                                                                          mem_19 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h13 == _T_158) begin
                                                                            mem_19 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h13 == _T_153) begin
                                                                              mem_19 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h13 == _T_308) begin
              mem_19 <= _GEN_31;
            end else begin
              if (6'h13 == _T_303) begin
                mem_19 <= _GEN_30;
              end else begin
                if (6'h13 == _T_298) begin
                  mem_19 <= _GEN_29;
                end else begin
                  if (6'h13 == _T_293) begin
                    mem_19 <= _GEN_28;
                  end else begin
                    if (6'h13 == _T_288) begin
                      mem_19 <= _GEN_27;
                    end else begin
                      if (6'h13 == _T_283) begin
                        mem_19 <= _GEN_26;
                      end else begin
                        if (6'h13 == _T_278) begin
                          mem_19 <= _GEN_25;
                        end else begin
                          if (6'h13 == _T_273) begin
                            mem_19 <= _GEN_24;
                          end else begin
                            if (6'h13 == _T_268) begin
                              mem_19 <= _GEN_23;
                            end else begin
                              if (6'h13 == _T_263) begin
                                mem_19 <= _GEN_22;
                              end else begin
                                if (6'h13 == _T_258) begin
                                  mem_19 <= _GEN_21;
                                end else begin
                                  if (6'h13 == _T_253) begin
                                    mem_19 <= _GEN_20;
                                  end else begin
                                    if (6'h13 == _T_248) begin
                                      mem_19 <= _GEN_19;
                                    end else begin
                                      if (6'h13 == _T_243) begin
                                        mem_19 <= _GEN_18;
                                      end else begin
                                        if (6'h13 == _T_238) begin
                                          mem_19 <= _GEN_17;
                                        end else begin
                                          if (6'h13 == _T_233) begin
                                            mem_19 <= _GEN_16;
                                          end else begin
                                            if (6'h13 == _T_228) begin
                                              mem_19 <= _GEN_15;
                                            end else begin
                                              if (6'h13 == _T_223) begin
                                                mem_19 <= _GEN_14;
                                              end else begin
                                                if (6'h13 == _T_218) begin
                                                  mem_19 <= _GEN_13;
                                                end else begin
                                                  if (6'h13 == _T_213) begin
                                                    mem_19 <= _GEN_12;
                                                  end else begin
                                                    if (6'h13 == _T_208) begin
                                                      mem_19 <= _GEN_11;
                                                    end else begin
                                                      if (6'h13 == _T_203) begin
                                                        mem_19 <= _GEN_10;
                                                      end else begin
                                                        if (6'h13 == _T_198) begin
                                                          mem_19 <= _GEN_9;
                                                        end else begin
                                                          if (6'h13 == _T_193) begin
                                                            mem_19 <= _GEN_8;
                                                          end else begin
                                                            if (6'h13 == _T_188) begin
                                                              mem_19 <= _GEN_7;
                                                            end else begin
                                                              if (6'h13 == _T_183) begin
                                                                mem_19 <= _GEN_6;
                                                              end else begin
                                                                if (6'h13 == _T_178) begin
                                                                  mem_19 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h13 == _T_173) begin
                                                                    mem_19 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h13 == _T_168) begin
                                                                      mem_19 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h13 == _T_163) begin
                                                                        mem_19 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h13 == _T_158) begin
                                                                          mem_19 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h13 == _T_153) begin
                                                                            mem_19 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h13 == _T_308) begin
            mem_19 <= _GEN_31;
          end else begin
            if (6'h13 == _T_303) begin
              mem_19 <= _GEN_30;
            end else begin
              if (6'h13 == _T_298) begin
                mem_19 <= _GEN_29;
              end else begin
                if (6'h13 == _T_293) begin
                  mem_19 <= _GEN_28;
                end else begin
                  if (6'h13 == _T_288) begin
                    mem_19 <= _GEN_27;
                  end else begin
                    if (6'h13 == _T_283) begin
                      mem_19 <= _GEN_26;
                    end else begin
                      if (6'h13 == _T_278) begin
                        mem_19 <= _GEN_25;
                      end else begin
                        if (6'h13 == _T_273) begin
                          mem_19 <= _GEN_24;
                        end else begin
                          if (6'h13 == _T_268) begin
                            mem_19 <= _GEN_23;
                          end else begin
                            if (6'h13 == _T_263) begin
                              mem_19 <= _GEN_22;
                            end else begin
                              if (6'h13 == _T_258) begin
                                mem_19 <= _GEN_21;
                              end else begin
                                if (6'h13 == _T_253) begin
                                  mem_19 <= _GEN_20;
                                end else begin
                                  if (6'h13 == _T_248) begin
                                    mem_19 <= _GEN_19;
                                  end else begin
                                    if (6'h13 == _T_243) begin
                                      mem_19 <= _GEN_18;
                                    end else begin
                                      if (6'h13 == _T_238) begin
                                        mem_19 <= _GEN_17;
                                      end else begin
                                        if (6'h13 == _T_233) begin
                                          mem_19 <= _GEN_16;
                                        end else begin
                                          if (6'h13 == _T_228) begin
                                            mem_19 <= _GEN_15;
                                          end else begin
                                            if (6'h13 == _T_223) begin
                                              mem_19 <= _GEN_14;
                                            end else begin
                                              if (6'h13 == _T_218) begin
                                                mem_19 <= _GEN_13;
                                              end else begin
                                                if (6'h13 == _T_213) begin
                                                  mem_19 <= _GEN_12;
                                                end else begin
                                                  if (6'h13 == _T_208) begin
                                                    mem_19 <= _GEN_11;
                                                  end else begin
                                                    if (6'h13 == _T_203) begin
                                                      mem_19 <= _GEN_10;
                                                    end else begin
                                                      if (6'h13 == _T_198) begin
                                                        mem_19 <= _GEN_9;
                                                      end else begin
                                                        if (6'h13 == _T_193) begin
                                                          mem_19 <= _GEN_8;
                                                        end else begin
                                                          if (6'h13 == _T_188) begin
                                                            mem_19 <= _GEN_7;
                                                          end else begin
                                                            if (6'h13 == _T_183) begin
                                                              mem_19 <= _GEN_6;
                                                            end else begin
                                                              if (6'h13 == _T_178) begin
                                                                mem_19 <= _GEN_5;
                                                              end else begin
                                                                if (6'h13 == _T_173) begin
                                                                  mem_19 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h13 == _T_168) begin
                                                                    mem_19 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h13 == _T_163) begin
                                                                      mem_19 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h13 == _T_158) begin
                                                                        mem_19 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h13 == _T_153) begin
                                                                          mem_19 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h13 == _T_308) begin
          mem_19 <= _GEN_31;
        end else begin
          if (6'h13 == _T_303) begin
            mem_19 <= _GEN_30;
          end else begin
            if (6'h13 == _T_298) begin
              mem_19 <= _GEN_29;
            end else begin
              if (6'h13 == _T_293) begin
                mem_19 <= _GEN_28;
              end else begin
                if (6'h13 == _T_288) begin
                  mem_19 <= _GEN_27;
                end else begin
                  if (6'h13 == _T_283) begin
                    mem_19 <= _GEN_26;
                  end else begin
                    if (6'h13 == _T_278) begin
                      mem_19 <= _GEN_25;
                    end else begin
                      if (6'h13 == _T_273) begin
                        mem_19 <= _GEN_24;
                      end else begin
                        if (6'h13 == _T_268) begin
                          mem_19 <= _GEN_23;
                        end else begin
                          if (6'h13 == _T_263) begin
                            mem_19 <= _GEN_22;
                          end else begin
                            if (6'h13 == _T_258) begin
                              mem_19 <= _GEN_21;
                            end else begin
                              if (6'h13 == _T_253) begin
                                mem_19 <= _GEN_20;
                              end else begin
                                if (6'h13 == _T_248) begin
                                  mem_19 <= _GEN_19;
                                end else begin
                                  if (6'h13 == _T_243) begin
                                    mem_19 <= _GEN_18;
                                  end else begin
                                    if (6'h13 == _T_238) begin
                                      mem_19 <= _GEN_17;
                                    end else begin
                                      if (6'h13 == _T_233) begin
                                        mem_19 <= _GEN_16;
                                      end else begin
                                        if (6'h13 == _T_228) begin
                                          mem_19 <= _GEN_15;
                                        end else begin
                                          if (6'h13 == _T_223) begin
                                            mem_19 <= _GEN_14;
                                          end else begin
                                            if (6'h13 == _T_218) begin
                                              mem_19 <= _GEN_13;
                                            end else begin
                                              if (6'h13 == _T_213) begin
                                                mem_19 <= _GEN_12;
                                              end else begin
                                                if (6'h13 == _T_208) begin
                                                  mem_19 <= _GEN_11;
                                                end else begin
                                                  if (6'h13 == _T_203) begin
                                                    mem_19 <= _GEN_10;
                                                  end else begin
                                                    if (6'h13 == _T_198) begin
                                                      mem_19 <= _GEN_9;
                                                    end else begin
                                                      if (6'h13 == _T_193) begin
                                                        mem_19 <= _GEN_8;
                                                      end else begin
                                                        if (6'h13 == _T_188) begin
                                                          mem_19 <= _GEN_7;
                                                        end else begin
                                                          if (6'h13 == _T_183) begin
                                                            mem_19 <= _GEN_6;
                                                          end else begin
                                                            if (6'h13 == _T_178) begin
                                                              mem_19 <= _GEN_5;
                                                            end else begin
                                                              if (6'h13 == _T_173) begin
                                                                mem_19 <= _GEN_4;
                                                              end else begin
                                                                if (6'h13 == _T_168) begin
                                                                  mem_19 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h13 == _T_163) begin
                                                                    mem_19 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h13 == _T_158) begin
                                                                      mem_19 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h13 == _T_153) begin
                                                                        mem_19 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h14 == wPos) begin
            mem_20 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h14 == _T_308) begin
                mem_20 <= _GEN_31;
              end else begin
                if (6'h14 == _T_303) begin
                  mem_20 <= _GEN_30;
                end else begin
                  if (6'h14 == _T_298) begin
                    mem_20 <= _GEN_29;
                  end else begin
                    if (6'h14 == _T_293) begin
                      mem_20 <= _GEN_28;
                    end else begin
                      if (6'h14 == _T_288) begin
                        mem_20 <= _GEN_27;
                      end else begin
                        if (6'h14 == _T_283) begin
                          mem_20 <= _GEN_26;
                        end else begin
                          if (6'h14 == _T_278) begin
                            mem_20 <= _GEN_25;
                          end else begin
                            if (6'h14 == _T_273) begin
                              mem_20 <= _GEN_24;
                            end else begin
                              if (6'h14 == _T_268) begin
                                mem_20 <= _GEN_23;
                              end else begin
                                if (6'h14 == _T_263) begin
                                  mem_20 <= _GEN_22;
                                end else begin
                                  if (6'h14 == _T_258) begin
                                    mem_20 <= _GEN_21;
                                  end else begin
                                    if (6'h14 == _T_253) begin
                                      mem_20 <= _GEN_20;
                                    end else begin
                                      if (6'h14 == _T_248) begin
                                        mem_20 <= _GEN_19;
                                      end else begin
                                        if (6'h14 == _T_243) begin
                                          mem_20 <= _GEN_18;
                                        end else begin
                                          if (6'h14 == _T_238) begin
                                            mem_20 <= _GEN_17;
                                          end else begin
                                            if (6'h14 == _T_233) begin
                                              mem_20 <= _GEN_16;
                                            end else begin
                                              if (6'h14 == _T_228) begin
                                                mem_20 <= _GEN_15;
                                              end else begin
                                                if (6'h14 == _T_223) begin
                                                  mem_20 <= _GEN_14;
                                                end else begin
                                                  if (6'h14 == _T_218) begin
                                                    mem_20 <= _GEN_13;
                                                  end else begin
                                                    if (6'h14 == _T_213) begin
                                                      mem_20 <= _GEN_12;
                                                    end else begin
                                                      if (6'h14 == _T_208) begin
                                                        mem_20 <= _GEN_11;
                                                      end else begin
                                                        if (6'h14 == _T_203) begin
                                                          mem_20 <= _GEN_10;
                                                        end else begin
                                                          if (6'h14 == _T_198) begin
                                                            mem_20 <= _GEN_9;
                                                          end else begin
                                                            if (6'h14 == _T_193) begin
                                                              mem_20 <= _GEN_8;
                                                            end else begin
                                                              if (6'h14 == _T_188) begin
                                                                mem_20 <= _GEN_7;
                                                              end else begin
                                                                if (6'h14 == _T_183) begin
                                                                  mem_20 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h14 == _T_178) begin
                                                                    mem_20 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h14 == _T_173) begin
                                                                      mem_20 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h14 == _T_168) begin
                                                                        mem_20 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h14 == _T_163) begin
                                                                          mem_20 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h14 == _T_158) begin
                                                                            mem_20 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h14 == _T_153) begin
                                                                              mem_20 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h14 == _T_308) begin
              mem_20 <= _GEN_31;
            end else begin
              if (6'h14 == _T_303) begin
                mem_20 <= _GEN_30;
              end else begin
                if (6'h14 == _T_298) begin
                  mem_20 <= _GEN_29;
                end else begin
                  if (6'h14 == _T_293) begin
                    mem_20 <= _GEN_28;
                  end else begin
                    if (6'h14 == _T_288) begin
                      mem_20 <= _GEN_27;
                    end else begin
                      if (6'h14 == _T_283) begin
                        mem_20 <= _GEN_26;
                      end else begin
                        if (6'h14 == _T_278) begin
                          mem_20 <= _GEN_25;
                        end else begin
                          if (6'h14 == _T_273) begin
                            mem_20 <= _GEN_24;
                          end else begin
                            if (6'h14 == _T_268) begin
                              mem_20 <= _GEN_23;
                            end else begin
                              if (6'h14 == _T_263) begin
                                mem_20 <= _GEN_22;
                              end else begin
                                if (6'h14 == _T_258) begin
                                  mem_20 <= _GEN_21;
                                end else begin
                                  if (6'h14 == _T_253) begin
                                    mem_20 <= _GEN_20;
                                  end else begin
                                    if (6'h14 == _T_248) begin
                                      mem_20 <= _GEN_19;
                                    end else begin
                                      if (6'h14 == _T_243) begin
                                        mem_20 <= _GEN_18;
                                      end else begin
                                        if (6'h14 == _T_238) begin
                                          mem_20 <= _GEN_17;
                                        end else begin
                                          if (6'h14 == _T_233) begin
                                            mem_20 <= _GEN_16;
                                          end else begin
                                            if (6'h14 == _T_228) begin
                                              mem_20 <= _GEN_15;
                                            end else begin
                                              if (6'h14 == _T_223) begin
                                                mem_20 <= _GEN_14;
                                              end else begin
                                                if (6'h14 == _T_218) begin
                                                  mem_20 <= _GEN_13;
                                                end else begin
                                                  if (6'h14 == _T_213) begin
                                                    mem_20 <= _GEN_12;
                                                  end else begin
                                                    if (6'h14 == _T_208) begin
                                                      mem_20 <= _GEN_11;
                                                    end else begin
                                                      if (6'h14 == _T_203) begin
                                                        mem_20 <= _GEN_10;
                                                      end else begin
                                                        if (6'h14 == _T_198) begin
                                                          mem_20 <= _GEN_9;
                                                        end else begin
                                                          if (6'h14 == _T_193) begin
                                                            mem_20 <= _GEN_8;
                                                          end else begin
                                                            if (6'h14 == _T_188) begin
                                                              mem_20 <= _GEN_7;
                                                            end else begin
                                                              if (6'h14 == _T_183) begin
                                                                mem_20 <= _GEN_6;
                                                              end else begin
                                                                if (6'h14 == _T_178) begin
                                                                  mem_20 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h14 == _T_173) begin
                                                                    mem_20 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h14 == _T_168) begin
                                                                      mem_20 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h14 == _T_163) begin
                                                                        mem_20 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h14 == _T_158) begin
                                                                          mem_20 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h14 == _T_153) begin
                                                                            mem_20 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h14 == _T_308) begin
            mem_20 <= _GEN_31;
          end else begin
            if (6'h14 == _T_303) begin
              mem_20 <= _GEN_30;
            end else begin
              if (6'h14 == _T_298) begin
                mem_20 <= _GEN_29;
              end else begin
                if (6'h14 == _T_293) begin
                  mem_20 <= _GEN_28;
                end else begin
                  if (6'h14 == _T_288) begin
                    mem_20 <= _GEN_27;
                  end else begin
                    if (6'h14 == _T_283) begin
                      mem_20 <= _GEN_26;
                    end else begin
                      if (6'h14 == _T_278) begin
                        mem_20 <= _GEN_25;
                      end else begin
                        if (6'h14 == _T_273) begin
                          mem_20 <= _GEN_24;
                        end else begin
                          if (6'h14 == _T_268) begin
                            mem_20 <= _GEN_23;
                          end else begin
                            if (6'h14 == _T_263) begin
                              mem_20 <= _GEN_22;
                            end else begin
                              if (6'h14 == _T_258) begin
                                mem_20 <= _GEN_21;
                              end else begin
                                if (6'h14 == _T_253) begin
                                  mem_20 <= _GEN_20;
                                end else begin
                                  if (6'h14 == _T_248) begin
                                    mem_20 <= _GEN_19;
                                  end else begin
                                    if (6'h14 == _T_243) begin
                                      mem_20 <= _GEN_18;
                                    end else begin
                                      if (6'h14 == _T_238) begin
                                        mem_20 <= _GEN_17;
                                      end else begin
                                        if (6'h14 == _T_233) begin
                                          mem_20 <= _GEN_16;
                                        end else begin
                                          if (6'h14 == _T_228) begin
                                            mem_20 <= _GEN_15;
                                          end else begin
                                            if (6'h14 == _T_223) begin
                                              mem_20 <= _GEN_14;
                                            end else begin
                                              if (6'h14 == _T_218) begin
                                                mem_20 <= _GEN_13;
                                              end else begin
                                                if (6'h14 == _T_213) begin
                                                  mem_20 <= _GEN_12;
                                                end else begin
                                                  if (6'h14 == _T_208) begin
                                                    mem_20 <= _GEN_11;
                                                  end else begin
                                                    if (6'h14 == _T_203) begin
                                                      mem_20 <= _GEN_10;
                                                    end else begin
                                                      if (6'h14 == _T_198) begin
                                                        mem_20 <= _GEN_9;
                                                      end else begin
                                                        if (6'h14 == _T_193) begin
                                                          mem_20 <= _GEN_8;
                                                        end else begin
                                                          if (6'h14 == _T_188) begin
                                                            mem_20 <= _GEN_7;
                                                          end else begin
                                                            if (6'h14 == _T_183) begin
                                                              mem_20 <= _GEN_6;
                                                            end else begin
                                                              if (6'h14 == _T_178) begin
                                                                mem_20 <= _GEN_5;
                                                              end else begin
                                                                if (6'h14 == _T_173) begin
                                                                  mem_20 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h14 == _T_168) begin
                                                                    mem_20 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h14 == _T_163) begin
                                                                      mem_20 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h14 == _T_158) begin
                                                                        mem_20 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h14 == _T_153) begin
                                                                          mem_20 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h14 == _T_308) begin
          mem_20 <= _GEN_31;
        end else begin
          if (6'h14 == _T_303) begin
            mem_20 <= _GEN_30;
          end else begin
            if (6'h14 == _T_298) begin
              mem_20 <= _GEN_29;
            end else begin
              if (6'h14 == _T_293) begin
                mem_20 <= _GEN_28;
              end else begin
                if (6'h14 == _T_288) begin
                  mem_20 <= _GEN_27;
                end else begin
                  if (6'h14 == _T_283) begin
                    mem_20 <= _GEN_26;
                  end else begin
                    if (6'h14 == _T_278) begin
                      mem_20 <= _GEN_25;
                    end else begin
                      if (6'h14 == _T_273) begin
                        mem_20 <= _GEN_24;
                      end else begin
                        if (6'h14 == _T_268) begin
                          mem_20 <= _GEN_23;
                        end else begin
                          if (6'h14 == _T_263) begin
                            mem_20 <= _GEN_22;
                          end else begin
                            if (6'h14 == _T_258) begin
                              mem_20 <= _GEN_21;
                            end else begin
                              if (6'h14 == _T_253) begin
                                mem_20 <= _GEN_20;
                              end else begin
                                if (6'h14 == _T_248) begin
                                  mem_20 <= _GEN_19;
                                end else begin
                                  if (6'h14 == _T_243) begin
                                    mem_20 <= _GEN_18;
                                  end else begin
                                    if (6'h14 == _T_238) begin
                                      mem_20 <= _GEN_17;
                                    end else begin
                                      if (6'h14 == _T_233) begin
                                        mem_20 <= _GEN_16;
                                      end else begin
                                        if (6'h14 == _T_228) begin
                                          mem_20 <= _GEN_15;
                                        end else begin
                                          if (6'h14 == _T_223) begin
                                            mem_20 <= _GEN_14;
                                          end else begin
                                            if (6'h14 == _T_218) begin
                                              mem_20 <= _GEN_13;
                                            end else begin
                                              if (6'h14 == _T_213) begin
                                                mem_20 <= _GEN_12;
                                              end else begin
                                                if (6'h14 == _T_208) begin
                                                  mem_20 <= _GEN_11;
                                                end else begin
                                                  if (6'h14 == _T_203) begin
                                                    mem_20 <= _GEN_10;
                                                  end else begin
                                                    if (6'h14 == _T_198) begin
                                                      mem_20 <= _GEN_9;
                                                    end else begin
                                                      if (6'h14 == _T_193) begin
                                                        mem_20 <= _GEN_8;
                                                      end else begin
                                                        if (6'h14 == _T_188) begin
                                                          mem_20 <= _GEN_7;
                                                        end else begin
                                                          if (6'h14 == _T_183) begin
                                                            mem_20 <= _GEN_6;
                                                          end else begin
                                                            if (6'h14 == _T_178) begin
                                                              mem_20 <= _GEN_5;
                                                            end else begin
                                                              if (6'h14 == _T_173) begin
                                                                mem_20 <= _GEN_4;
                                                              end else begin
                                                                if (6'h14 == _T_168) begin
                                                                  mem_20 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h14 == _T_163) begin
                                                                    mem_20 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h14 == _T_158) begin
                                                                      mem_20 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h14 == _T_153) begin
                                                                        mem_20 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h15 == wPos) begin
            mem_21 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h15 == _T_308) begin
                mem_21 <= _GEN_31;
              end else begin
                if (6'h15 == _T_303) begin
                  mem_21 <= _GEN_30;
                end else begin
                  if (6'h15 == _T_298) begin
                    mem_21 <= _GEN_29;
                  end else begin
                    if (6'h15 == _T_293) begin
                      mem_21 <= _GEN_28;
                    end else begin
                      if (6'h15 == _T_288) begin
                        mem_21 <= _GEN_27;
                      end else begin
                        if (6'h15 == _T_283) begin
                          mem_21 <= _GEN_26;
                        end else begin
                          if (6'h15 == _T_278) begin
                            mem_21 <= _GEN_25;
                          end else begin
                            if (6'h15 == _T_273) begin
                              mem_21 <= _GEN_24;
                            end else begin
                              if (6'h15 == _T_268) begin
                                mem_21 <= _GEN_23;
                              end else begin
                                if (6'h15 == _T_263) begin
                                  mem_21 <= _GEN_22;
                                end else begin
                                  if (6'h15 == _T_258) begin
                                    mem_21 <= _GEN_21;
                                  end else begin
                                    if (6'h15 == _T_253) begin
                                      mem_21 <= _GEN_20;
                                    end else begin
                                      if (6'h15 == _T_248) begin
                                        mem_21 <= _GEN_19;
                                      end else begin
                                        if (6'h15 == _T_243) begin
                                          mem_21 <= _GEN_18;
                                        end else begin
                                          if (6'h15 == _T_238) begin
                                            mem_21 <= _GEN_17;
                                          end else begin
                                            if (6'h15 == _T_233) begin
                                              mem_21 <= _GEN_16;
                                            end else begin
                                              if (6'h15 == _T_228) begin
                                                mem_21 <= _GEN_15;
                                              end else begin
                                                if (6'h15 == _T_223) begin
                                                  mem_21 <= _GEN_14;
                                                end else begin
                                                  if (6'h15 == _T_218) begin
                                                    mem_21 <= _GEN_13;
                                                  end else begin
                                                    if (6'h15 == _T_213) begin
                                                      mem_21 <= _GEN_12;
                                                    end else begin
                                                      if (6'h15 == _T_208) begin
                                                        mem_21 <= _GEN_11;
                                                      end else begin
                                                        if (6'h15 == _T_203) begin
                                                          mem_21 <= _GEN_10;
                                                        end else begin
                                                          if (6'h15 == _T_198) begin
                                                            mem_21 <= _GEN_9;
                                                          end else begin
                                                            if (6'h15 == _T_193) begin
                                                              mem_21 <= _GEN_8;
                                                            end else begin
                                                              if (6'h15 == _T_188) begin
                                                                mem_21 <= _GEN_7;
                                                              end else begin
                                                                if (6'h15 == _T_183) begin
                                                                  mem_21 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h15 == _T_178) begin
                                                                    mem_21 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h15 == _T_173) begin
                                                                      mem_21 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h15 == _T_168) begin
                                                                        mem_21 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h15 == _T_163) begin
                                                                          mem_21 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h15 == _T_158) begin
                                                                            mem_21 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h15 == _T_153) begin
                                                                              mem_21 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h15 == _T_308) begin
              mem_21 <= _GEN_31;
            end else begin
              if (6'h15 == _T_303) begin
                mem_21 <= _GEN_30;
              end else begin
                if (6'h15 == _T_298) begin
                  mem_21 <= _GEN_29;
                end else begin
                  if (6'h15 == _T_293) begin
                    mem_21 <= _GEN_28;
                  end else begin
                    if (6'h15 == _T_288) begin
                      mem_21 <= _GEN_27;
                    end else begin
                      if (6'h15 == _T_283) begin
                        mem_21 <= _GEN_26;
                      end else begin
                        if (6'h15 == _T_278) begin
                          mem_21 <= _GEN_25;
                        end else begin
                          if (6'h15 == _T_273) begin
                            mem_21 <= _GEN_24;
                          end else begin
                            if (6'h15 == _T_268) begin
                              mem_21 <= _GEN_23;
                            end else begin
                              if (6'h15 == _T_263) begin
                                mem_21 <= _GEN_22;
                              end else begin
                                if (6'h15 == _T_258) begin
                                  mem_21 <= _GEN_21;
                                end else begin
                                  if (6'h15 == _T_253) begin
                                    mem_21 <= _GEN_20;
                                  end else begin
                                    if (6'h15 == _T_248) begin
                                      mem_21 <= _GEN_19;
                                    end else begin
                                      if (6'h15 == _T_243) begin
                                        mem_21 <= _GEN_18;
                                      end else begin
                                        if (6'h15 == _T_238) begin
                                          mem_21 <= _GEN_17;
                                        end else begin
                                          if (6'h15 == _T_233) begin
                                            mem_21 <= _GEN_16;
                                          end else begin
                                            if (6'h15 == _T_228) begin
                                              mem_21 <= _GEN_15;
                                            end else begin
                                              if (6'h15 == _T_223) begin
                                                mem_21 <= _GEN_14;
                                              end else begin
                                                if (6'h15 == _T_218) begin
                                                  mem_21 <= _GEN_13;
                                                end else begin
                                                  if (6'h15 == _T_213) begin
                                                    mem_21 <= _GEN_12;
                                                  end else begin
                                                    if (6'h15 == _T_208) begin
                                                      mem_21 <= _GEN_11;
                                                    end else begin
                                                      if (6'h15 == _T_203) begin
                                                        mem_21 <= _GEN_10;
                                                      end else begin
                                                        if (6'h15 == _T_198) begin
                                                          mem_21 <= _GEN_9;
                                                        end else begin
                                                          if (6'h15 == _T_193) begin
                                                            mem_21 <= _GEN_8;
                                                          end else begin
                                                            if (6'h15 == _T_188) begin
                                                              mem_21 <= _GEN_7;
                                                            end else begin
                                                              if (6'h15 == _T_183) begin
                                                                mem_21 <= _GEN_6;
                                                              end else begin
                                                                if (6'h15 == _T_178) begin
                                                                  mem_21 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h15 == _T_173) begin
                                                                    mem_21 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h15 == _T_168) begin
                                                                      mem_21 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h15 == _T_163) begin
                                                                        mem_21 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h15 == _T_158) begin
                                                                          mem_21 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h15 == _T_153) begin
                                                                            mem_21 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h15 == _T_308) begin
            mem_21 <= _GEN_31;
          end else begin
            if (6'h15 == _T_303) begin
              mem_21 <= _GEN_30;
            end else begin
              if (6'h15 == _T_298) begin
                mem_21 <= _GEN_29;
              end else begin
                if (6'h15 == _T_293) begin
                  mem_21 <= _GEN_28;
                end else begin
                  if (6'h15 == _T_288) begin
                    mem_21 <= _GEN_27;
                  end else begin
                    if (6'h15 == _T_283) begin
                      mem_21 <= _GEN_26;
                    end else begin
                      if (6'h15 == _T_278) begin
                        mem_21 <= _GEN_25;
                      end else begin
                        if (6'h15 == _T_273) begin
                          mem_21 <= _GEN_24;
                        end else begin
                          if (6'h15 == _T_268) begin
                            mem_21 <= _GEN_23;
                          end else begin
                            if (6'h15 == _T_263) begin
                              mem_21 <= _GEN_22;
                            end else begin
                              if (6'h15 == _T_258) begin
                                mem_21 <= _GEN_21;
                              end else begin
                                if (6'h15 == _T_253) begin
                                  mem_21 <= _GEN_20;
                                end else begin
                                  if (6'h15 == _T_248) begin
                                    mem_21 <= _GEN_19;
                                  end else begin
                                    if (6'h15 == _T_243) begin
                                      mem_21 <= _GEN_18;
                                    end else begin
                                      if (6'h15 == _T_238) begin
                                        mem_21 <= _GEN_17;
                                      end else begin
                                        if (6'h15 == _T_233) begin
                                          mem_21 <= _GEN_16;
                                        end else begin
                                          if (6'h15 == _T_228) begin
                                            mem_21 <= _GEN_15;
                                          end else begin
                                            if (6'h15 == _T_223) begin
                                              mem_21 <= _GEN_14;
                                            end else begin
                                              if (6'h15 == _T_218) begin
                                                mem_21 <= _GEN_13;
                                              end else begin
                                                if (6'h15 == _T_213) begin
                                                  mem_21 <= _GEN_12;
                                                end else begin
                                                  if (6'h15 == _T_208) begin
                                                    mem_21 <= _GEN_11;
                                                  end else begin
                                                    if (6'h15 == _T_203) begin
                                                      mem_21 <= _GEN_10;
                                                    end else begin
                                                      if (6'h15 == _T_198) begin
                                                        mem_21 <= _GEN_9;
                                                      end else begin
                                                        if (6'h15 == _T_193) begin
                                                          mem_21 <= _GEN_8;
                                                        end else begin
                                                          if (6'h15 == _T_188) begin
                                                            mem_21 <= _GEN_7;
                                                          end else begin
                                                            if (6'h15 == _T_183) begin
                                                              mem_21 <= _GEN_6;
                                                            end else begin
                                                              if (6'h15 == _T_178) begin
                                                                mem_21 <= _GEN_5;
                                                              end else begin
                                                                if (6'h15 == _T_173) begin
                                                                  mem_21 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h15 == _T_168) begin
                                                                    mem_21 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h15 == _T_163) begin
                                                                      mem_21 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h15 == _T_158) begin
                                                                        mem_21 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h15 == _T_153) begin
                                                                          mem_21 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h15 == _T_308) begin
          mem_21 <= _GEN_31;
        end else begin
          if (6'h15 == _T_303) begin
            mem_21 <= _GEN_30;
          end else begin
            if (6'h15 == _T_298) begin
              mem_21 <= _GEN_29;
            end else begin
              if (6'h15 == _T_293) begin
                mem_21 <= _GEN_28;
              end else begin
                if (6'h15 == _T_288) begin
                  mem_21 <= _GEN_27;
                end else begin
                  if (6'h15 == _T_283) begin
                    mem_21 <= _GEN_26;
                  end else begin
                    if (6'h15 == _T_278) begin
                      mem_21 <= _GEN_25;
                    end else begin
                      if (6'h15 == _T_273) begin
                        mem_21 <= _GEN_24;
                      end else begin
                        if (6'h15 == _T_268) begin
                          mem_21 <= _GEN_23;
                        end else begin
                          if (6'h15 == _T_263) begin
                            mem_21 <= _GEN_22;
                          end else begin
                            if (6'h15 == _T_258) begin
                              mem_21 <= _GEN_21;
                            end else begin
                              if (6'h15 == _T_253) begin
                                mem_21 <= _GEN_20;
                              end else begin
                                if (6'h15 == _T_248) begin
                                  mem_21 <= _GEN_19;
                                end else begin
                                  if (6'h15 == _T_243) begin
                                    mem_21 <= _GEN_18;
                                  end else begin
                                    if (6'h15 == _T_238) begin
                                      mem_21 <= _GEN_17;
                                    end else begin
                                      if (6'h15 == _T_233) begin
                                        mem_21 <= _GEN_16;
                                      end else begin
                                        if (6'h15 == _T_228) begin
                                          mem_21 <= _GEN_15;
                                        end else begin
                                          if (6'h15 == _T_223) begin
                                            mem_21 <= _GEN_14;
                                          end else begin
                                            if (6'h15 == _T_218) begin
                                              mem_21 <= _GEN_13;
                                            end else begin
                                              if (6'h15 == _T_213) begin
                                                mem_21 <= _GEN_12;
                                              end else begin
                                                if (6'h15 == _T_208) begin
                                                  mem_21 <= _GEN_11;
                                                end else begin
                                                  if (6'h15 == _T_203) begin
                                                    mem_21 <= _GEN_10;
                                                  end else begin
                                                    if (6'h15 == _T_198) begin
                                                      mem_21 <= _GEN_9;
                                                    end else begin
                                                      if (6'h15 == _T_193) begin
                                                        mem_21 <= _GEN_8;
                                                      end else begin
                                                        if (6'h15 == _T_188) begin
                                                          mem_21 <= _GEN_7;
                                                        end else begin
                                                          if (6'h15 == _T_183) begin
                                                            mem_21 <= _GEN_6;
                                                          end else begin
                                                            if (6'h15 == _T_178) begin
                                                              mem_21 <= _GEN_5;
                                                            end else begin
                                                              if (6'h15 == _T_173) begin
                                                                mem_21 <= _GEN_4;
                                                              end else begin
                                                                if (6'h15 == _T_168) begin
                                                                  mem_21 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h15 == _T_163) begin
                                                                    mem_21 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h15 == _T_158) begin
                                                                      mem_21 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h15 == _T_153) begin
                                                                        mem_21 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h16 == wPos) begin
            mem_22 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h16 == _T_308) begin
                mem_22 <= _GEN_31;
              end else begin
                if (6'h16 == _T_303) begin
                  mem_22 <= _GEN_30;
                end else begin
                  if (6'h16 == _T_298) begin
                    mem_22 <= _GEN_29;
                  end else begin
                    if (6'h16 == _T_293) begin
                      mem_22 <= _GEN_28;
                    end else begin
                      if (6'h16 == _T_288) begin
                        mem_22 <= _GEN_27;
                      end else begin
                        if (6'h16 == _T_283) begin
                          mem_22 <= _GEN_26;
                        end else begin
                          if (6'h16 == _T_278) begin
                            mem_22 <= _GEN_25;
                          end else begin
                            if (6'h16 == _T_273) begin
                              mem_22 <= _GEN_24;
                            end else begin
                              if (6'h16 == _T_268) begin
                                mem_22 <= _GEN_23;
                              end else begin
                                if (6'h16 == _T_263) begin
                                  mem_22 <= _GEN_22;
                                end else begin
                                  if (6'h16 == _T_258) begin
                                    mem_22 <= _GEN_21;
                                  end else begin
                                    if (6'h16 == _T_253) begin
                                      mem_22 <= _GEN_20;
                                    end else begin
                                      if (6'h16 == _T_248) begin
                                        mem_22 <= _GEN_19;
                                      end else begin
                                        if (6'h16 == _T_243) begin
                                          mem_22 <= _GEN_18;
                                        end else begin
                                          if (6'h16 == _T_238) begin
                                            mem_22 <= _GEN_17;
                                          end else begin
                                            if (6'h16 == _T_233) begin
                                              mem_22 <= _GEN_16;
                                            end else begin
                                              if (6'h16 == _T_228) begin
                                                mem_22 <= _GEN_15;
                                              end else begin
                                                if (6'h16 == _T_223) begin
                                                  mem_22 <= _GEN_14;
                                                end else begin
                                                  if (6'h16 == _T_218) begin
                                                    mem_22 <= _GEN_13;
                                                  end else begin
                                                    if (6'h16 == _T_213) begin
                                                      mem_22 <= _GEN_12;
                                                    end else begin
                                                      if (6'h16 == _T_208) begin
                                                        mem_22 <= _GEN_11;
                                                      end else begin
                                                        if (6'h16 == _T_203) begin
                                                          mem_22 <= _GEN_10;
                                                        end else begin
                                                          if (6'h16 == _T_198) begin
                                                            mem_22 <= _GEN_9;
                                                          end else begin
                                                            if (6'h16 == _T_193) begin
                                                              mem_22 <= _GEN_8;
                                                            end else begin
                                                              if (6'h16 == _T_188) begin
                                                                mem_22 <= _GEN_7;
                                                              end else begin
                                                                if (6'h16 == _T_183) begin
                                                                  mem_22 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h16 == _T_178) begin
                                                                    mem_22 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h16 == _T_173) begin
                                                                      mem_22 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h16 == _T_168) begin
                                                                        mem_22 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h16 == _T_163) begin
                                                                          mem_22 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h16 == _T_158) begin
                                                                            mem_22 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h16 == _T_153) begin
                                                                              mem_22 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h16 == _T_308) begin
              mem_22 <= _GEN_31;
            end else begin
              if (6'h16 == _T_303) begin
                mem_22 <= _GEN_30;
              end else begin
                if (6'h16 == _T_298) begin
                  mem_22 <= _GEN_29;
                end else begin
                  if (6'h16 == _T_293) begin
                    mem_22 <= _GEN_28;
                  end else begin
                    if (6'h16 == _T_288) begin
                      mem_22 <= _GEN_27;
                    end else begin
                      if (6'h16 == _T_283) begin
                        mem_22 <= _GEN_26;
                      end else begin
                        if (6'h16 == _T_278) begin
                          mem_22 <= _GEN_25;
                        end else begin
                          if (6'h16 == _T_273) begin
                            mem_22 <= _GEN_24;
                          end else begin
                            if (6'h16 == _T_268) begin
                              mem_22 <= _GEN_23;
                            end else begin
                              if (6'h16 == _T_263) begin
                                mem_22 <= _GEN_22;
                              end else begin
                                if (6'h16 == _T_258) begin
                                  mem_22 <= _GEN_21;
                                end else begin
                                  if (6'h16 == _T_253) begin
                                    mem_22 <= _GEN_20;
                                  end else begin
                                    if (6'h16 == _T_248) begin
                                      mem_22 <= _GEN_19;
                                    end else begin
                                      if (6'h16 == _T_243) begin
                                        mem_22 <= _GEN_18;
                                      end else begin
                                        if (6'h16 == _T_238) begin
                                          mem_22 <= _GEN_17;
                                        end else begin
                                          if (6'h16 == _T_233) begin
                                            mem_22 <= _GEN_16;
                                          end else begin
                                            if (6'h16 == _T_228) begin
                                              mem_22 <= _GEN_15;
                                            end else begin
                                              if (6'h16 == _T_223) begin
                                                mem_22 <= _GEN_14;
                                              end else begin
                                                if (6'h16 == _T_218) begin
                                                  mem_22 <= _GEN_13;
                                                end else begin
                                                  if (6'h16 == _T_213) begin
                                                    mem_22 <= _GEN_12;
                                                  end else begin
                                                    if (6'h16 == _T_208) begin
                                                      mem_22 <= _GEN_11;
                                                    end else begin
                                                      if (6'h16 == _T_203) begin
                                                        mem_22 <= _GEN_10;
                                                      end else begin
                                                        if (6'h16 == _T_198) begin
                                                          mem_22 <= _GEN_9;
                                                        end else begin
                                                          if (6'h16 == _T_193) begin
                                                            mem_22 <= _GEN_8;
                                                          end else begin
                                                            if (6'h16 == _T_188) begin
                                                              mem_22 <= _GEN_7;
                                                            end else begin
                                                              if (6'h16 == _T_183) begin
                                                                mem_22 <= _GEN_6;
                                                              end else begin
                                                                if (6'h16 == _T_178) begin
                                                                  mem_22 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h16 == _T_173) begin
                                                                    mem_22 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h16 == _T_168) begin
                                                                      mem_22 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h16 == _T_163) begin
                                                                        mem_22 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h16 == _T_158) begin
                                                                          mem_22 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h16 == _T_153) begin
                                                                            mem_22 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h16 == _T_308) begin
            mem_22 <= _GEN_31;
          end else begin
            if (6'h16 == _T_303) begin
              mem_22 <= _GEN_30;
            end else begin
              if (6'h16 == _T_298) begin
                mem_22 <= _GEN_29;
              end else begin
                if (6'h16 == _T_293) begin
                  mem_22 <= _GEN_28;
                end else begin
                  if (6'h16 == _T_288) begin
                    mem_22 <= _GEN_27;
                  end else begin
                    if (6'h16 == _T_283) begin
                      mem_22 <= _GEN_26;
                    end else begin
                      if (6'h16 == _T_278) begin
                        mem_22 <= _GEN_25;
                      end else begin
                        if (6'h16 == _T_273) begin
                          mem_22 <= _GEN_24;
                        end else begin
                          if (6'h16 == _T_268) begin
                            mem_22 <= _GEN_23;
                          end else begin
                            if (6'h16 == _T_263) begin
                              mem_22 <= _GEN_22;
                            end else begin
                              if (6'h16 == _T_258) begin
                                mem_22 <= _GEN_21;
                              end else begin
                                if (6'h16 == _T_253) begin
                                  mem_22 <= _GEN_20;
                                end else begin
                                  if (6'h16 == _T_248) begin
                                    mem_22 <= _GEN_19;
                                  end else begin
                                    if (6'h16 == _T_243) begin
                                      mem_22 <= _GEN_18;
                                    end else begin
                                      if (6'h16 == _T_238) begin
                                        mem_22 <= _GEN_17;
                                      end else begin
                                        if (6'h16 == _T_233) begin
                                          mem_22 <= _GEN_16;
                                        end else begin
                                          if (6'h16 == _T_228) begin
                                            mem_22 <= _GEN_15;
                                          end else begin
                                            if (6'h16 == _T_223) begin
                                              mem_22 <= _GEN_14;
                                            end else begin
                                              if (6'h16 == _T_218) begin
                                                mem_22 <= _GEN_13;
                                              end else begin
                                                if (6'h16 == _T_213) begin
                                                  mem_22 <= _GEN_12;
                                                end else begin
                                                  if (6'h16 == _T_208) begin
                                                    mem_22 <= _GEN_11;
                                                  end else begin
                                                    if (6'h16 == _T_203) begin
                                                      mem_22 <= _GEN_10;
                                                    end else begin
                                                      if (6'h16 == _T_198) begin
                                                        mem_22 <= _GEN_9;
                                                      end else begin
                                                        if (6'h16 == _T_193) begin
                                                          mem_22 <= _GEN_8;
                                                        end else begin
                                                          if (6'h16 == _T_188) begin
                                                            mem_22 <= _GEN_7;
                                                          end else begin
                                                            if (6'h16 == _T_183) begin
                                                              mem_22 <= _GEN_6;
                                                            end else begin
                                                              if (6'h16 == _T_178) begin
                                                                mem_22 <= _GEN_5;
                                                              end else begin
                                                                if (6'h16 == _T_173) begin
                                                                  mem_22 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h16 == _T_168) begin
                                                                    mem_22 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h16 == _T_163) begin
                                                                      mem_22 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h16 == _T_158) begin
                                                                        mem_22 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h16 == _T_153) begin
                                                                          mem_22 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h16 == _T_308) begin
          mem_22 <= _GEN_31;
        end else begin
          if (6'h16 == _T_303) begin
            mem_22 <= _GEN_30;
          end else begin
            if (6'h16 == _T_298) begin
              mem_22 <= _GEN_29;
            end else begin
              if (6'h16 == _T_293) begin
                mem_22 <= _GEN_28;
              end else begin
                if (6'h16 == _T_288) begin
                  mem_22 <= _GEN_27;
                end else begin
                  if (6'h16 == _T_283) begin
                    mem_22 <= _GEN_26;
                  end else begin
                    if (6'h16 == _T_278) begin
                      mem_22 <= _GEN_25;
                    end else begin
                      if (6'h16 == _T_273) begin
                        mem_22 <= _GEN_24;
                      end else begin
                        if (6'h16 == _T_268) begin
                          mem_22 <= _GEN_23;
                        end else begin
                          if (6'h16 == _T_263) begin
                            mem_22 <= _GEN_22;
                          end else begin
                            if (6'h16 == _T_258) begin
                              mem_22 <= _GEN_21;
                            end else begin
                              if (6'h16 == _T_253) begin
                                mem_22 <= _GEN_20;
                              end else begin
                                if (6'h16 == _T_248) begin
                                  mem_22 <= _GEN_19;
                                end else begin
                                  if (6'h16 == _T_243) begin
                                    mem_22 <= _GEN_18;
                                  end else begin
                                    if (6'h16 == _T_238) begin
                                      mem_22 <= _GEN_17;
                                    end else begin
                                      if (6'h16 == _T_233) begin
                                        mem_22 <= _GEN_16;
                                      end else begin
                                        if (6'h16 == _T_228) begin
                                          mem_22 <= _GEN_15;
                                        end else begin
                                          if (6'h16 == _T_223) begin
                                            mem_22 <= _GEN_14;
                                          end else begin
                                            if (6'h16 == _T_218) begin
                                              mem_22 <= _GEN_13;
                                            end else begin
                                              if (6'h16 == _T_213) begin
                                                mem_22 <= _GEN_12;
                                              end else begin
                                                if (6'h16 == _T_208) begin
                                                  mem_22 <= _GEN_11;
                                                end else begin
                                                  if (6'h16 == _T_203) begin
                                                    mem_22 <= _GEN_10;
                                                  end else begin
                                                    if (6'h16 == _T_198) begin
                                                      mem_22 <= _GEN_9;
                                                    end else begin
                                                      if (6'h16 == _T_193) begin
                                                        mem_22 <= _GEN_8;
                                                      end else begin
                                                        if (6'h16 == _T_188) begin
                                                          mem_22 <= _GEN_7;
                                                        end else begin
                                                          if (6'h16 == _T_183) begin
                                                            mem_22 <= _GEN_6;
                                                          end else begin
                                                            if (6'h16 == _T_178) begin
                                                              mem_22 <= _GEN_5;
                                                            end else begin
                                                              if (6'h16 == _T_173) begin
                                                                mem_22 <= _GEN_4;
                                                              end else begin
                                                                if (6'h16 == _T_168) begin
                                                                  mem_22 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h16 == _T_163) begin
                                                                    mem_22 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h16 == _T_158) begin
                                                                      mem_22 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h16 == _T_153) begin
                                                                        mem_22 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h17 == wPos) begin
            mem_23 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h17 == _T_308) begin
                mem_23 <= _GEN_31;
              end else begin
                if (6'h17 == _T_303) begin
                  mem_23 <= _GEN_30;
                end else begin
                  if (6'h17 == _T_298) begin
                    mem_23 <= _GEN_29;
                  end else begin
                    if (6'h17 == _T_293) begin
                      mem_23 <= _GEN_28;
                    end else begin
                      if (6'h17 == _T_288) begin
                        mem_23 <= _GEN_27;
                      end else begin
                        if (6'h17 == _T_283) begin
                          mem_23 <= _GEN_26;
                        end else begin
                          if (6'h17 == _T_278) begin
                            mem_23 <= _GEN_25;
                          end else begin
                            if (6'h17 == _T_273) begin
                              mem_23 <= _GEN_24;
                            end else begin
                              if (6'h17 == _T_268) begin
                                mem_23 <= _GEN_23;
                              end else begin
                                if (6'h17 == _T_263) begin
                                  mem_23 <= _GEN_22;
                                end else begin
                                  if (6'h17 == _T_258) begin
                                    mem_23 <= _GEN_21;
                                  end else begin
                                    if (6'h17 == _T_253) begin
                                      mem_23 <= _GEN_20;
                                    end else begin
                                      if (6'h17 == _T_248) begin
                                        mem_23 <= _GEN_19;
                                      end else begin
                                        if (6'h17 == _T_243) begin
                                          mem_23 <= _GEN_18;
                                        end else begin
                                          if (6'h17 == _T_238) begin
                                            mem_23 <= _GEN_17;
                                          end else begin
                                            if (6'h17 == _T_233) begin
                                              mem_23 <= _GEN_16;
                                            end else begin
                                              if (6'h17 == _T_228) begin
                                                mem_23 <= _GEN_15;
                                              end else begin
                                                if (6'h17 == _T_223) begin
                                                  mem_23 <= _GEN_14;
                                                end else begin
                                                  if (6'h17 == _T_218) begin
                                                    mem_23 <= _GEN_13;
                                                  end else begin
                                                    if (6'h17 == _T_213) begin
                                                      mem_23 <= _GEN_12;
                                                    end else begin
                                                      if (6'h17 == _T_208) begin
                                                        mem_23 <= _GEN_11;
                                                      end else begin
                                                        if (6'h17 == _T_203) begin
                                                          mem_23 <= _GEN_10;
                                                        end else begin
                                                          if (6'h17 == _T_198) begin
                                                            mem_23 <= _GEN_9;
                                                          end else begin
                                                            if (6'h17 == _T_193) begin
                                                              mem_23 <= _GEN_8;
                                                            end else begin
                                                              if (6'h17 == _T_188) begin
                                                                mem_23 <= _GEN_7;
                                                              end else begin
                                                                if (6'h17 == _T_183) begin
                                                                  mem_23 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h17 == _T_178) begin
                                                                    mem_23 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h17 == _T_173) begin
                                                                      mem_23 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h17 == _T_168) begin
                                                                        mem_23 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h17 == _T_163) begin
                                                                          mem_23 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h17 == _T_158) begin
                                                                            mem_23 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h17 == _T_153) begin
                                                                              mem_23 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h17 == _T_308) begin
              mem_23 <= _GEN_31;
            end else begin
              if (6'h17 == _T_303) begin
                mem_23 <= _GEN_30;
              end else begin
                if (6'h17 == _T_298) begin
                  mem_23 <= _GEN_29;
                end else begin
                  if (6'h17 == _T_293) begin
                    mem_23 <= _GEN_28;
                  end else begin
                    if (6'h17 == _T_288) begin
                      mem_23 <= _GEN_27;
                    end else begin
                      if (6'h17 == _T_283) begin
                        mem_23 <= _GEN_26;
                      end else begin
                        if (6'h17 == _T_278) begin
                          mem_23 <= _GEN_25;
                        end else begin
                          if (6'h17 == _T_273) begin
                            mem_23 <= _GEN_24;
                          end else begin
                            if (6'h17 == _T_268) begin
                              mem_23 <= _GEN_23;
                            end else begin
                              if (6'h17 == _T_263) begin
                                mem_23 <= _GEN_22;
                              end else begin
                                if (6'h17 == _T_258) begin
                                  mem_23 <= _GEN_21;
                                end else begin
                                  if (6'h17 == _T_253) begin
                                    mem_23 <= _GEN_20;
                                  end else begin
                                    if (6'h17 == _T_248) begin
                                      mem_23 <= _GEN_19;
                                    end else begin
                                      if (6'h17 == _T_243) begin
                                        mem_23 <= _GEN_18;
                                      end else begin
                                        if (6'h17 == _T_238) begin
                                          mem_23 <= _GEN_17;
                                        end else begin
                                          if (6'h17 == _T_233) begin
                                            mem_23 <= _GEN_16;
                                          end else begin
                                            if (6'h17 == _T_228) begin
                                              mem_23 <= _GEN_15;
                                            end else begin
                                              if (6'h17 == _T_223) begin
                                                mem_23 <= _GEN_14;
                                              end else begin
                                                if (6'h17 == _T_218) begin
                                                  mem_23 <= _GEN_13;
                                                end else begin
                                                  if (6'h17 == _T_213) begin
                                                    mem_23 <= _GEN_12;
                                                  end else begin
                                                    if (6'h17 == _T_208) begin
                                                      mem_23 <= _GEN_11;
                                                    end else begin
                                                      if (6'h17 == _T_203) begin
                                                        mem_23 <= _GEN_10;
                                                      end else begin
                                                        if (6'h17 == _T_198) begin
                                                          mem_23 <= _GEN_9;
                                                        end else begin
                                                          if (6'h17 == _T_193) begin
                                                            mem_23 <= _GEN_8;
                                                          end else begin
                                                            if (6'h17 == _T_188) begin
                                                              mem_23 <= _GEN_7;
                                                            end else begin
                                                              if (6'h17 == _T_183) begin
                                                                mem_23 <= _GEN_6;
                                                              end else begin
                                                                if (6'h17 == _T_178) begin
                                                                  mem_23 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h17 == _T_173) begin
                                                                    mem_23 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h17 == _T_168) begin
                                                                      mem_23 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h17 == _T_163) begin
                                                                        mem_23 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h17 == _T_158) begin
                                                                          mem_23 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h17 == _T_153) begin
                                                                            mem_23 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h17 == _T_308) begin
            mem_23 <= _GEN_31;
          end else begin
            if (6'h17 == _T_303) begin
              mem_23 <= _GEN_30;
            end else begin
              if (6'h17 == _T_298) begin
                mem_23 <= _GEN_29;
              end else begin
                if (6'h17 == _T_293) begin
                  mem_23 <= _GEN_28;
                end else begin
                  if (6'h17 == _T_288) begin
                    mem_23 <= _GEN_27;
                  end else begin
                    if (6'h17 == _T_283) begin
                      mem_23 <= _GEN_26;
                    end else begin
                      if (6'h17 == _T_278) begin
                        mem_23 <= _GEN_25;
                      end else begin
                        if (6'h17 == _T_273) begin
                          mem_23 <= _GEN_24;
                        end else begin
                          if (6'h17 == _T_268) begin
                            mem_23 <= _GEN_23;
                          end else begin
                            if (6'h17 == _T_263) begin
                              mem_23 <= _GEN_22;
                            end else begin
                              if (6'h17 == _T_258) begin
                                mem_23 <= _GEN_21;
                              end else begin
                                if (6'h17 == _T_253) begin
                                  mem_23 <= _GEN_20;
                                end else begin
                                  if (6'h17 == _T_248) begin
                                    mem_23 <= _GEN_19;
                                  end else begin
                                    if (6'h17 == _T_243) begin
                                      mem_23 <= _GEN_18;
                                    end else begin
                                      if (6'h17 == _T_238) begin
                                        mem_23 <= _GEN_17;
                                      end else begin
                                        if (6'h17 == _T_233) begin
                                          mem_23 <= _GEN_16;
                                        end else begin
                                          if (6'h17 == _T_228) begin
                                            mem_23 <= _GEN_15;
                                          end else begin
                                            if (6'h17 == _T_223) begin
                                              mem_23 <= _GEN_14;
                                            end else begin
                                              if (6'h17 == _T_218) begin
                                                mem_23 <= _GEN_13;
                                              end else begin
                                                if (6'h17 == _T_213) begin
                                                  mem_23 <= _GEN_12;
                                                end else begin
                                                  if (6'h17 == _T_208) begin
                                                    mem_23 <= _GEN_11;
                                                  end else begin
                                                    if (6'h17 == _T_203) begin
                                                      mem_23 <= _GEN_10;
                                                    end else begin
                                                      if (6'h17 == _T_198) begin
                                                        mem_23 <= _GEN_9;
                                                      end else begin
                                                        if (6'h17 == _T_193) begin
                                                          mem_23 <= _GEN_8;
                                                        end else begin
                                                          if (6'h17 == _T_188) begin
                                                            mem_23 <= _GEN_7;
                                                          end else begin
                                                            if (6'h17 == _T_183) begin
                                                              mem_23 <= _GEN_6;
                                                            end else begin
                                                              if (6'h17 == _T_178) begin
                                                                mem_23 <= _GEN_5;
                                                              end else begin
                                                                if (6'h17 == _T_173) begin
                                                                  mem_23 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h17 == _T_168) begin
                                                                    mem_23 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h17 == _T_163) begin
                                                                      mem_23 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h17 == _T_158) begin
                                                                        mem_23 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h17 == _T_153) begin
                                                                          mem_23 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h17 == _T_308) begin
          mem_23 <= _GEN_31;
        end else begin
          if (6'h17 == _T_303) begin
            mem_23 <= _GEN_30;
          end else begin
            if (6'h17 == _T_298) begin
              mem_23 <= _GEN_29;
            end else begin
              if (6'h17 == _T_293) begin
                mem_23 <= _GEN_28;
              end else begin
                if (6'h17 == _T_288) begin
                  mem_23 <= _GEN_27;
                end else begin
                  if (6'h17 == _T_283) begin
                    mem_23 <= _GEN_26;
                  end else begin
                    if (6'h17 == _T_278) begin
                      mem_23 <= _GEN_25;
                    end else begin
                      if (6'h17 == _T_273) begin
                        mem_23 <= _GEN_24;
                      end else begin
                        if (6'h17 == _T_268) begin
                          mem_23 <= _GEN_23;
                        end else begin
                          if (6'h17 == _T_263) begin
                            mem_23 <= _GEN_22;
                          end else begin
                            if (6'h17 == _T_258) begin
                              mem_23 <= _GEN_21;
                            end else begin
                              if (6'h17 == _T_253) begin
                                mem_23 <= _GEN_20;
                              end else begin
                                if (6'h17 == _T_248) begin
                                  mem_23 <= _GEN_19;
                                end else begin
                                  if (6'h17 == _T_243) begin
                                    mem_23 <= _GEN_18;
                                  end else begin
                                    if (6'h17 == _T_238) begin
                                      mem_23 <= _GEN_17;
                                    end else begin
                                      if (6'h17 == _T_233) begin
                                        mem_23 <= _GEN_16;
                                      end else begin
                                        if (6'h17 == _T_228) begin
                                          mem_23 <= _GEN_15;
                                        end else begin
                                          if (6'h17 == _T_223) begin
                                            mem_23 <= _GEN_14;
                                          end else begin
                                            if (6'h17 == _T_218) begin
                                              mem_23 <= _GEN_13;
                                            end else begin
                                              if (6'h17 == _T_213) begin
                                                mem_23 <= _GEN_12;
                                              end else begin
                                                if (6'h17 == _T_208) begin
                                                  mem_23 <= _GEN_11;
                                                end else begin
                                                  if (6'h17 == _T_203) begin
                                                    mem_23 <= _GEN_10;
                                                  end else begin
                                                    if (6'h17 == _T_198) begin
                                                      mem_23 <= _GEN_9;
                                                    end else begin
                                                      if (6'h17 == _T_193) begin
                                                        mem_23 <= _GEN_8;
                                                      end else begin
                                                        if (6'h17 == _T_188) begin
                                                          mem_23 <= _GEN_7;
                                                        end else begin
                                                          if (6'h17 == _T_183) begin
                                                            mem_23 <= _GEN_6;
                                                          end else begin
                                                            if (6'h17 == _T_178) begin
                                                              mem_23 <= _GEN_5;
                                                            end else begin
                                                              if (6'h17 == _T_173) begin
                                                                mem_23 <= _GEN_4;
                                                              end else begin
                                                                if (6'h17 == _T_168) begin
                                                                  mem_23 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h17 == _T_163) begin
                                                                    mem_23 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h17 == _T_158) begin
                                                                      mem_23 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h17 == _T_153) begin
                                                                        mem_23 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h18 == wPos) begin
            mem_24 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h18 == _T_308) begin
                mem_24 <= _GEN_31;
              end else begin
                if (6'h18 == _T_303) begin
                  mem_24 <= _GEN_30;
                end else begin
                  if (6'h18 == _T_298) begin
                    mem_24 <= _GEN_29;
                  end else begin
                    if (6'h18 == _T_293) begin
                      mem_24 <= _GEN_28;
                    end else begin
                      if (6'h18 == _T_288) begin
                        mem_24 <= _GEN_27;
                      end else begin
                        if (6'h18 == _T_283) begin
                          mem_24 <= _GEN_26;
                        end else begin
                          if (6'h18 == _T_278) begin
                            mem_24 <= _GEN_25;
                          end else begin
                            if (6'h18 == _T_273) begin
                              mem_24 <= _GEN_24;
                            end else begin
                              if (6'h18 == _T_268) begin
                                mem_24 <= _GEN_23;
                              end else begin
                                if (6'h18 == _T_263) begin
                                  mem_24 <= _GEN_22;
                                end else begin
                                  if (6'h18 == _T_258) begin
                                    mem_24 <= _GEN_21;
                                  end else begin
                                    if (6'h18 == _T_253) begin
                                      mem_24 <= _GEN_20;
                                    end else begin
                                      if (6'h18 == _T_248) begin
                                        mem_24 <= _GEN_19;
                                      end else begin
                                        if (6'h18 == _T_243) begin
                                          mem_24 <= _GEN_18;
                                        end else begin
                                          if (6'h18 == _T_238) begin
                                            mem_24 <= _GEN_17;
                                          end else begin
                                            if (6'h18 == _T_233) begin
                                              mem_24 <= _GEN_16;
                                            end else begin
                                              if (6'h18 == _T_228) begin
                                                mem_24 <= _GEN_15;
                                              end else begin
                                                if (6'h18 == _T_223) begin
                                                  mem_24 <= _GEN_14;
                                                end else begin
                                                  if (6'h18 == _T_218) begin
                                                    mem_24 <= _GEN_13;
                                                  end else begin
                                                    if (6'h18 == _T_213) begin
                                                      mem_24 <= _GEN_12;
                                                    end else begin
                                                      if (6'h18 == _T_208) begin
                                                        mem_24 <= _GEN_11;
                                                      end else begin
                                                        if (6'h18 == _T_203) begin
                                                          mem_24 <= _GEN_10;
                                                        end else begin
                                                          if (6'h18 == _T_198) begin
                                                            mem_24 <= _GEN_9;
                                                          end else begin
                                                            if (6'h18 == _T_193) begin
                                                              mem_24 <= _GEN_8;
                                                            end else begin
                                                              if (6'h18 == _T_188) begin
                                                                mem_24 <= _GEN_7;
                                                              end else begin
                                                                if (6'h18 == _T_183) begin
                                                                  mem_24 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h18 == _T_178) begin
                                                                    mem_24 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h18 == _T_173) begin
                                                                      mem_24 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h18 == _T_168) begin
                                                                        mem_24 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h18 == _T_163) begin
                                                                          mem_24 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h18 == _T_158) begin
                                                                            mem_24 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h18 == _T_153) begin
                                                                              mem_24 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h18 == _T_308) begin
              mem_24 <= _GEN_31;
            end else begin
              if (6'h18 == _T_303) begin
                mem_24 <= _GEN_30;
              end else begin
                if (6'h18 == _T_298) begin
                  mem_24 <= _GEN_29;
                end else begin
                  if (6'h18 == _T_293) begin
                    mem_24 <= _GEN_28;
                  end else begin
                    if (6'h18 == _T_288) begin
                      mem_24 <= _GEN_27;
                    end else begin
                      if (6'h18 == _T_283) begin
                        mem_24 <= _GEN_26;
                      end else begin
                        if (6'h18 == _T_278) begin
                          mem_24 <= _GEN_25;
                        end else begin
                          if (6'h18 == _T_273) begin
                            mem_24 <= _GEN_24;
                          end else begin
                            if (6'h18 == _T_268) begin
                              mem_24 <= _GEN_23;
                            end else begin
                              if (6'h18 == _T_263) begin
                                mem_24 <= _GEN_22;
                              end else begin
                                if (6'h18 == _T_258) begin
                                  mem_24 <= _GEN_21;
                                end else begin
                                  if (6'h18 == _T_253) begin
                                    mem_24 <= _GEN_20;
                                  end else begin
                                    if (6'h18 == _T_248) begin
                                      mem_24 <= _GEN_19;
                                    end else begin
                                      if (6'h18 == _T_243) begin
                                        mem_24 <= _GEN_18;
                                      end else begin
                                        if (6'h18 == _T_238) begin
                                          mem_24 <= _GEN_17;
                                        end else begin
                                          if (6'h18 == _T_233) begin
                                            mem_24 <= _GEN_16;
                                          end else begin
                                            if (6'h18 == _T_228) begin
                                              mem_24 <= _GEN_15;
                                            end else begin
                                              if (6'h18 == _T_223) begin
                                                mem_24 <= _GEN_14;
                                              end else begin
                                                if (6'h18 == _T_218) begin
                                                  mem_24 <= _GEN_13;
                                                end else begin
                                                  if (6'h18 == _T_213) begin
                                                    mem_24 <= _GEN_12;
                                                  end else begin
                                                    if (6'h18 == _T_208) begin
                                                      mem_24 <= _GEN_11;
                                                    end else begin
                                                      if (6'h18 == _T_203) begin
                                                        mem_24 <= _GEN_10;
                                                      end else begin
                                                        if (6'h18 == _T_198) begin
                                                          mem_24 <= _GEN_9;
                                                        end else begin
                                                          if (6'h18 == _T_193) begin
                                                            mem_24 <= _GEN_8;
                                                          end else begin
                                                            if (6'h18 == _T_188) begin
                                                              mem_24 <= _GEN_7;
                                                            end else begin
                                                              if (6'h18 == _T_183) begin
                                                                mem_24 <= _GEN_6;
                                                              end else begin
                                                                if (6'h18 == _T_178) begin
                                                                  mem_24 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h18 == _T_173) begin
                                                                    mem_24 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h18 == _T_168) begin
                                                                      mem_24 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h18 == _T_163) begin
                                                                        mem_24 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h18 == _T_158) begin
                                                                          mem_24 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h18 == _T_153) begin
                                                                            mem_24 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h18 == _T_308) begin
            mem_24 <= _GEN_31;
          end else begin
            if (6'h18 == _T_303) begin
              mem_24 <= _GEN_30;
            end else begin
              if (6'h18 == _T_298) begin
                mem_24 <= _GEN_29;
              end else begin
                if (6'h18 == _T_293) begin
                  mem_24 <= _GEN_28;
                end else begin
                  if (6'h18 == _T_288) begin
                    mem_24 <= _GEN_27;
                  end else begin
                    if (6'h18 == _T_283) begin
                      mem_24 <= _GEN_26;
                    end else begin
                      if (6'h18 == _T_278) begin
                        mem_24 <= _GEN_25;
                      end else begin
                        if (6'h18 == _T_273) begin
                          mem_24 <= _GEN_24;
                        end else begin
                          if (6'h18 == _T_268) begin
                            mem_24 <= _GEN_23;
                          end else begin
                            if (6'h18 == _T_263) begin
                              mem_24 <= _GEN_22;
                            end else begin
                              if (6'h18 == _T_258) begin
                                mem_24 <= _GEN_21;
                              end else begin
                                if (6'h18 == _T_253) begin
                                  mem_24 <= _GEN_20;
                                end else begin
                                  if (6'h18 == _T_248) begin
                                    mem_24 <= _GEN_19;
                                  end else begin
                                    if (6'h18 == _T_243) begin
                                      mem_24 <= _GEN_18;
                                    end else begin
                                      if (6'h18 == _T_238) begin
                                        mem_24 <= _GEN_17;
                                      end else begin
                                        if (6'h18 == _T_233) begin
                                          mem_24 <= _GEN_16;
                                        end else begin
                                          if (6'h18 == _T_228) begin
                                            mem_24 <= _GEN_15;
                                          end else begin
                                            if (6'h18 == _T_223) begin
                                              mem_24 <= _GEN_14;
                                            end else begin
                                              if (6'h18 == _T_218) begin
                                                mem_24 <= _GEN_13;
                                              end else begin
                                                if (6'h18 == _T_213) begin
                                                  mem_24 <= _GEN_12;
                                                end else begin
                                                  if (6'h18 == _T_208) begin
                                                    mem_24 <= _GEN_11;
                                                  end else begin
                                                    if (6'h18 == _T_203) begin
                                                      mem_24 <= _GEN_10;
                                                    end else begin
                                                      if (6'h18 == _T_198) begin
                                                        mem_24 <= _GEN_9;
                                                      end else begin
                                                        if (6'h18 == _T_193) begin
                                                          mem_24 <= _GEN_8;
                                                        end else begin
                                                          if (6'h18 == _T_188) begin
                                                            mem_24 <= _GEN_7;
                                                          end else begin
                                                            if (6'h18 == _T_183) begin
                                                              mem_24 <= _GEN_6;
                                                            end else begin
                                                              if (6'h18 == _T_178) begin
                                                                mem_24 <= _GEN_5;
                                                              end else begin
                                                                if (6'h18 == _T_173) begin
                                                                  mem_24 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h18 == _T_168) begin
                                                                    mem_24 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h18 == _T_163) begin
                                                                      mem_24 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h18 == _T_158) begin
                                                                        mem_24 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h18 == _T_153) begin
                                                                          mem_24 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h18 == _T_308) begin
          mem_24 <= _GEN_31;
        end else begin
          if (6'h18 == _T_303) begin
            mem_24 <= _GEN_30;
          end else begin
            if (6'h18 == _T_298) begin
              mem_24 <= _GEN_29;
            end else begin
              if (6'h18 == _T_293) begin
                mem_24 <= _GEN_28;
              end else begin
                if (6'h18 == _T_288) begin
                  mem_24 <= _GEN_27;
                end else begin
                  if (6'h18 == _T_283) begin
                    mem_24 <= _GEN_26;
                  end else begin
                    if (6'h18 == _T_278) begin
                      mem_24 <= _GEN_25;
                    end else begin
                      if (6'h18 == _T_273) begin
                        mem_24 <= _GEN_24;
                      end else begin
                        if (6'h18 == _T_268) begin
                          mem_24 <= _GEN_23;
                        end else begin
                          if (6'h18 == _T_263) begin
                            mem_24 <= _GEN_22;
                          end else begin
                            if (6'h18 == _T_258) begin
                              mem_24 <= _GEN_21;
                            end else begin
                              if (6'h18 == _T_253) begin
                                mem_24 <= _GEN_20;
                              end else begin
                                if (6'h18 == _T_248) begin
                                  mem_24 <= _GEN_19;
                                end else begin
                                  if (6'h18 == _T_243) begin
                                    mem_24 <= _GEN_18;
                                  end else begin
                                    if (6'h18 == _T_238) begin
                                      mem_24 <= _GEN_17;
                                    end else begin
                                      if (6'h18 == _T_233) begin
                                        mem_24 <= _GEN_16;
                                      end else begin
                                        if (6'h18 == _T_228) begin
                                          mem_24 <= _GEN_15;
                                        end else begin
                                          if (6'h18 == _T_223) begin
                                            mem_24 <= _GEN_14;
                                          end else begin
                                            if (6'h18 == _T_218) begin
                                              mem_24 <= _GEN_13;
                                            end else begin
                                              if (6'h18 == _T_213) begin
                                                mem_24 <= _GEN_12;
                                              end else begin
                                                if (6'h18 == _T_208) begin
                                                  mem_24 <= _GEN_11;
                                                end else begin
                                                  if (6'h18 == _T_203) begin
                                                    mem_24 <= _GEN_10;
                                                  end else begin
                                                    if (6'h18 == _T_198) begin
                                                      mem_24 <= _GEN_9;
                                                    end else begin
                                                      if (6'h18 == _T_193) begin
                                                        mem_24 <= _GEN_8;
                                                      end else begin
                                                        if (6'h18 == _T_188) begin
                                                          mem_24 <= _GEN_7;
                                                        end else begin
                                                          if (6'h18 == _T_183) begin
                                                            mem_24 <= _GEN_6;
                                                          end else begin
                                                            if (6'h18 == _T_178) begin
                                                              mem_24 <= _GEN_5;
                                                            end else begin
                                                              if (6'h18 == _T_173) begin
                                                                mem_24 <= _GEN_4;
                                                              end else begin
                                                                if (6'h18 == _T_168) begin
                                                                  mem_24 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h18 == _T_163) begin
                                                                    mem_24 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h18 == _T_158) begin
                                                                      mem_24 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h18 == _T_153) begin
                                                                        mem_24 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h19 == wPos) begin
            mem_25 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h19 == _T_308) begin
                mem_25 <= _GEN_31;
              end else begin
                if (6'h19 == _T_303) begin
                  mem_25 <= _GEN_30;
                end else begin
                  if (6'h19 == _T_298) begin
                    mem_25 <= _GEN_29;
                  end else begin
                    if (6'h19 == _T_293) begin
                      mem_25 <= _GEN_28;
                    end else begin
                      if (6'h19 == _T_288) begin
                        mem_25 <= _GEN_27;
                      end else begin
                        if (6'h19 == _T_283) begin
                          mem_25 <= _GEN_26;
                        end else begin
                          if (6'h19 == _T_278) begin
                            mem_25 <= _GEN_25;
                          end else begin
                            if (6'h19 == _T_273) begin
                              mem_25 <= _GEN_24;
                            end else begin
                              if (6'h19 == _T_268) begin
                                mem_25 <= _GEN_23;
                              end else begin
                                if (6'h19 == _T_263) begin
                                  mem_25 <= _GEN_22;
                                end else begin
                                  if (6'h19 == _T_258) begin
                                    mem_25 <= _GEN_21;
                                  end else begin
                                    if (6'h19 == _T_253) begin
                                      mem_25 <= _GEN_20;
                                    end else begin
                                      if (6'h19 == _T_248) begin
                                        mem_25 <= _GEN_19;
                                      end else begin
                                        if (6'h19 == _T_243) begin
                                          mem_25 <= _GEN_18;
                                        end else begin
                                          if (6'h19 == _T_238) begin
                                            mem_25 <= _GEN_17;
                                          end else begin
                                            if (6'h19 == _T_233) begin
                                              mem_25 <= _GEN_16;
                                            end else begin
                                              if (6'h19 == _T_228) begin
                                                mem_25 <= _GEN_15;
                                              end else begin
                                                if (6'h19 == _T_223) begin
                                                  mem_25 <= _GEN_14;
                                                end else begin
                                                  if (6'h19 == _T_218) begin
                                                    mem_25 <= _GEN_13;
                                                  end else begin
                                                    if (6'h19 == _T_213) begin
                                                      mem_25 <= _GEN_12;
                                                    end else begin
                                                      if (6'h19 == _T_208) begin
                                                        mem_25 <= _GEN_11;
                                                      end else begin
                                                        if (6'h19 == _T_203) begin
                                                          mem_25 <= _GEN_10;
                                                        end else begin
                                                          if (6'h19 == _T_198) begin
                                                            mem_25 <= _GEN_9;
                                                          end else begin
                                                            if (6'h19 == _T_193) begin
                                                              mem_25 <= _GEN_8;
                                                            end else begin
                                                              if (6'h19 == _T_188) begin
                                                                mem_25 <= _GEN_7;
                                                              end else begin
                                                                if (6'h19 == _T_183) begin
                                                                  mem_25 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h19 == _T_178) begin
                                                                    mem_25 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h19 == _T_173) begin
                                                                      mem_25 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h19 == _T_168) begin
                                                                        mem_25 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h19 == _T_163) begin
                                                                          mem_25 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h19 == _T_158) begin
                                                                            mem_25 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h19 == _T_153) begin
                                                                              mem_25 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h19 == _T_308) begin
              mem_25 <= _GEN_31;
            end else begin
              if (6'h19 == _T_303) begin
                mem_25 <= _GEN_30;
              end else begin
                if (6'h19 == _T_298) begin
                  mem_25 <= _GEN_29;
                end else begin
                  if (6'h19 == _T_293) begin
                    mem_25 <= _GEN_28;
                  end else begin
                    if (6'h19 == _T_288) begin
                      mem_25 <= _GEN_27;
                    end else begin
                      if (6'h19 == _T_283) begin
                        mem_25 <= _GEN_26;
                      end else begin
                        if (6'h19 == _T_278) begin
                          mem_25 <= _GEN_25;
                        end else begin
                          if (6'h19 == _T_273) begin
                            mem_25 <= _GEN_24;
                          end else begin
                            if (6'h19 == _T_268) begin
                              mem_25 <= _GEN_23;
                            end else begin
                              if (6'h19 == _T_263) begin
                                mem_25 <= _GEN_22;
                              end else begin
                                if (6'h19 == _T_258) begin
                                  mem_25 <= _GEN_21;
                                end else begin
                                  if (6'h19 == _T_253) begin
                                    mem_25 <= _GEN_20;
                                  end else begin
                                    if (6'h19 == _T_248) begin
                                      mem_25 <= _GEN_19;
                                    end else begin
                                      if (6'h19 == _T_243) begin
                                        mem_25 <= _GEN_18;
                                      end else begin
                                        if (6'h19 == _T_238) begin
                                          mem_25 <= _GEN_17;
                                        end else begin
                                          if (6'h19 == _T_233) begin
                                            mem_25 <= _GEN_16;
                                          end else begin
                                            if (6'h19 == _T_228) begin
                                              mem_25 <= _GEN_15;
                                            end else begin
                                              if (6'h19 == _T_223) begin
                                                mem_25 <= _GEN_14;
                                              end else begin
                                                if (6'h19 == _T_218) begin
                                                  mem_25 <= _GEN_13;
                                                end else begin
                                                  if (6'h19 == _T_213) begin
                                                    mem_25 <= _GEN_12;
                                                  end else begin
                                                    if (6'h19 == _T_208) begin
                                                      mem_25 <= _GEN_11;
                                                    end else begin
                                                      if (6'h19 == _T_203) begin
                                                        mem_25 <= _GEN_10;
                                                      end else begin
                                                        if (6'h19 == _T_198) begin
                                                          mem_25 <= _GEN_9;
                                                        end else begin
                                                          if (6'h19 == _T_193) begin
                                                            mem_25 <= _GEN_8;
                                                          end else begin
                                                            if (6'h19 == _T_188) begin
                                                              mem_25 <= _GEN_7;
                                                            end else begin
                                                              if (6'h19 == _T_183) begin
                                                                mem_25 <= _GEN_6;
                                                              end else begin
                                                                if (6'h19 == _T_178) begin
                                                                  mem_25 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h19 == _T_173) begin
                                                                    mem_25 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h19 == _T_168) begin
                                                                      mem_25 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h19 == _T_163) begin
                                                                        mem_25 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h19 == _T_158) begin
                                                                          mem_25 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h19 == _T_153) begin
                                                                            mem_25 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h19 == _T_308) begin
            mem_25 <= _GEN_31;
          end else begin
            if (6'h19 == _T_303) begin
              mem_25 <= _GEN_30;
            end else begin
              if (6'h19 == _T_298) begin
                mem_25 <= _GEN_29;
              end else begin
                if (6'h19 == _T_293) begin
                  mem_25 <= _GEN_28;
                end else begin
                  if (6'h19 == _T_288) begin
                    mem_25 <= _GEN_27;
                  end else begin
                    if (6'h19 == _T_283) begin
                      mem_25 <= _GEN_26;
                    end else begin
                      if (6'h19 == _T_278) begin
                        mem_25 <= _GEN_25;
                      end else begin
                        if (6'h19 == _T_273) begin
                          mem_25 <= _GEN_24;
                        end else begin
                          if (6'h19 == _T_268) begin
                            mem_25 <= _GEN_23;
                          end else begin
                            if (6'h19 == _T_263) begin
                              mem_25 <= _GEN_22;
                            end else begin
                              if (6'h19 == _T_258) begin
                                mem_25 <= _GEN_21;
                              end else begin
                                if (6'h19 == _T_253) begin
                                  mem_25 <= _GEN_20;
                                end else begin
                                  if (6'h19 == _T_248) begin
                                    mem_25 <= _GEN_19;
                                  end else begin
                                    if (6'h19 == _T_243) begin
                                      mem_25 <= _GEN_18;
                                    end else begin
                                      if (6'h19 == _T_238) begin
                                        mem_25 <= _GEN_17;
                                      end else begin
                                        if (6'h19 == _T_233) begin
                                          mem_25 <= _GEN_16;
                                        end else begin
                                          if (6'h19 == _T_228) begin
                                            mem_25 <= _GEN_15;
                                          end else begin
                                            if (6'h19 == _T_223) begin
                                              mem_25 <= _GEN_14;
                                            end else begin
                                              if (6'h19 == _T_218) begin
                                                mem_25 <= _GEN_13;
                                              end else begin
                                                if (6'h19 == _T_213) begin
                                                  mem_25 <= _GEN_12;
                                                end else begin
                                                  if (6'h19 == _T_208) begin
                                                    mem_25 <= _GEN_11;
                                                  end else begin
                                                    if (6'h19 == _T_203) begin
                                                      mem_25 <= _GEN_10;
                                                    end else begin
                                                      if (6'h19 == _T_198) begin
                                                        mem_25 <= _GEN_9;
                                                      end else begin
                                                        if (6'h19 == _T_193) begin
                                                          mem_25 <= _GEN_8;
                                                        end else begin
                                                          if (6'h19 == _T_188) begin
                                                            mem_25 <= _GEN_7;
                                                          end else begin
                                                            if (6'h19 == _T_183) begin
                                                              mem_25 <= _GEN_6;
                                                            end else begin
                                                              if (6'h19 == _T_178) begin
                                                                mem_25 <= _GEN_5;
                                                              end else begin
                                                                if (6'h19 == _T_173) begin
                                                                  mem_25 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h19 == _T_168) begin
                                                                    mem_25 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h19 == _T_163) begin
                                                                      mem_25 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h19 == _T_158) begin
                                                                        mem_25 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h19 == _T_153) begin
                                                                          mem_25 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h19 == _T_308) begin
          mem_25 <= _GEN_31;
        end else begin
          if (6'h19 == _T_303) begin
            mem_25 <= _GEN_30;
          end else begin
            if (6'h19 == _T_298) begin
              mem_25 <= _GEN_29;
            end else begin
              if (6'h19 == _T_293) begin
                mem_25 <= _GEN_28;
              end else begin
                if (6'h19 == _T_288) begin
                  mem_25 <= _GEN_27;
                end else begin
                  if (6'h19 == _T_283) begin
                    mem_25 <= _GEN_26;
                  end else begin
                    if (6'h19 == _T_278) begin
                      mem_25 <= _GEN_25;
                    end else begin
                      if (6'h19 == _T_273) begin
                        mem_25 <= _GEN_24;
                      end else begin
                        if (6'h19 == _T_268) begin
                          mem_25 <= _GEN_23;
                        end else begin
                          if (6'h19 == _T_263) begin
                            mem_25 <= _GEN_22;
                          end else begin
                            if (6'h19 == _T_258) begin
                              mem_25 <= _GEN_21;
                            end else begin
                              if (6'h19 == _T_253) begin
                                mem_25 <= _GEN_20;
                              end else begin
                                if (6'h19 == _T_248) begin
                                  mem_25 <= _GEN_19;
                                end else begin
                                  if (6'h19 == _T_243) begin
                                    mem_25 <= _GEN_18;
                                  end else begin
                                    if (6'h19 == _T_238) begin
                                      mem_25 <= _GEN_17;
                                    end else begin
                                      if (6'h19 == _T_233) begin
                                        mem_25 <= _GEN_16;
                                      end else begin
                                        if (6'h19 == _T_228) begin
                                          mem_25 <= _GEN_15;
                                        end else begin
                                          if (6'h19 == _T_223) begin
                                            mem_25 <= _GEN_14;
                                          end else begin
                                            if (6'h19 == _T_218) begin
                                              mem_25 <= _GEN_13;
                                            end else begin
                                              if (6'h19 == _T_213) begin
                                                mem_25 <= _GEN_12;
                                              end else begin
                                                if (6'h19 == _T_208) begin
                                                  mem_25 <= _GEN_11;
                                                end else begin
                                                  if (6'h19 == _T_203) begin
                                                    mem_25 <= _GEN_10;
                                                  end else begin
                                                    if (6'h19 == _T_198) begin
                                                      mem_25 <= _GEN_9;
                                                    end else begin
                                                      if (6'h19 == _T_193) begin
                                                        mem_25 <= _GEN_8;
                                                      end else begin
                                                        if (6'h19 == _T_188) begin
                                                          mem_25 <= _GEN_7;
                                                        end else begin
                                                          if (6'h19 == _T_183) begin
                                                            mem_25 <= _GEN_6;
                                                          end else begin
                                                            if (6'h19 == _T_178) begin
                                                              mem_25 <= _GEN_5;
                                                            end else begin
                                                              if (6'h19 == _T_173) begin
                                                                mem_25 <= _GEN_4;
                                                              end else begin
                                                                if (6'h19 == _T_168) begin
                                                                  mem_25 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h19 == _T_163) begin
                                                                    mem_25 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h19 == _T_158) begin
                                                                      mem_25 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h19 == _T_153) begin
                                                                        mem_25 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h1a == wPos) begin
            mem_26 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h1a == _T_308) begin
                mem_26 <= _GEN_31;
              end else begin
                if (6'h1a == _T_303) begin
                  mem_26 <= _GEN_30;
                end else begin
                  if (6'h1a == _T_298) begin
                    mem_26 <= _GEN_29;
                  end else begin
                    if (6'h1a == _T_293) begin
                      mem_26 <= _GEN_28;
                    end else begin
                      if (6'h1a == _T_288) begin
                        mem_26 <= _GEN_27;
                      end else begin
                        if (6'h1a == _T_283) begin
                          mem_26 <= _GEN_26;
                        end else begin
                          if (6'h1a == _T_278) begin
                            mem_26 <= _GEN_25;
                          end else begin
                            if (6'h1a == _T_273) begin
                              mem_26 <= _GEN_24;
                            end else begin
                              if (6'h1a == _T_268) begin
                                mem_26 <= _GEN_23;
                              end else begin
                                if (6'h1a == _T_263) begin
                                  mem_26 <= _GEN_22;
                                end else begin
                                  if (6'h1a == _T_258) begin
                                    mem_26 <= _GEN_21;
                                  end else begin
                                    if (6'h1a == _T_253) begin
                                      mem_26 <= _GEN_20;
                                    end else begin
                                      if (6'h1a == _T_248) begin
                                        mem_26 <= _GEN_19;
                                      end else begin
                                        if (6'h1a == _T_243) begin
                                          mem_26 <= _GEN_18;
                                        end else begin
                                          if (6'h1a == _T_238) begin
                                            mem_26 <= _GEN_17;
                                          end else begin
                                            if (6'h1a == _T_233) begin
                                              mem_26 <= _GEN_16;
                                            end else begin
                                              if (6'h1a == _T_228) begin
                                                mem_26 <= _GEN_15;
                                              end else begin
                                                if (6'h1a == _T_223) begin
                                                  mem_26 <= _GEN_14;
                                                end else begin
                                                  if (6'h1a == _T_218) begin
                                                    mem_26 <= _GEN_13;
                                                  end else begin
                                                    if (6'h1a == _T_213) begin
                                                      mem_26 <= _GEN_12;
                                                    end else begin
                                                      if (6'h1a == _T_208) begin
                                                        mem_26 <= _GEN_11;
                                                      end else begin
                                                        if (6'h1a == _T_203) begin
                                                          mem_26 <= _GEN_10;
                                                        end else begin
                                                          if (6'h1a == _T_198) begin
                                                            mem_26 <= _GEN_9;
                                                          end else begin
                                                            if (6'h1a == _T_193) begin
                                                              mem_26 <= _GEN_8;
                                                            end else begin
                                                              if (6'h1a == _T_188) begin
                                                                mem_26 <= _GEN_7;
                                                              end else begin
                                                                if (6'h1a == _T_183) begin
                                                                  mem_26 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h1a == _T_178) begin
                                                                    mem_26 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h1a == _T_173) begin
                                                                      mem_26 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h1a == _T_168) begin
                                                                        mem_26 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h1a == _T_163) begin
                                                                          mem_26 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h1a == _T_158) begin
                                                                            mem_26 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h1a == _T_153) begin
                                                                              mem_26 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h1a == _T_308) begin
              mem_26 <= _GEN_31;
            end else begin
              if (6'h1a == _T_303) begin
                mem_26 <= _GEN_30;
              end else begin
                if (6'h1a == _T_298) begin
                  mem_26 <= _GEN_29;
                end else begin
                  if (6'h1a == _T_293) begin
                    mem_26 <= _GEN_28;
                  end else begin
                    if (6'h1a == _T_288) begin
                      mem_26 <= _GEN_27;
                    end else begin
                      if (6'h1a == _T_283) begin
                        mem_26 <= _GEN_26;
                      end else begin
                        if (6'h1a == _T_278) begin
                          mem_26 <= _GEN_25;
                        end else begin
                          if (6'h1a == _T_273) begin
                            mem_26 <= _GEN_24;
                          end else begin
                            if (6'h1a == _T_268) begin
                              mem_26 <= _GEN_23;
                            end else begin
                              if (6'h1a == _T_263) begin
                                mem_26 <= _GEN_22;
                              end else begin
                                if (6'h1a == _T_258) begin
                                  mem_26 <= _GEN_21;
                                end else begin
                                  if (6'h1a == _T_253) begin
                                    mem_26 <= _GEN_20;
                                  end else begin
                                    if (6'h1a == _T_248) begin
                                      mem_26 <= _GEN_19;
                                    end else begin
                                      if (6'h1a == _T_243) begin
                                        mem_26 <= _GEN_18;
                                      end else begin
                                        if (6'h1a == _T_238) begin
                                          mem_26 <= _GEN_17;
                                        end else begin
                                          if (6'h1a == _T_233) begin
                                            mem_26 <= _GEN_16;
                                          end else begin
                                            if (6'h1a == _T_228) begin
                                              mem_26 <= _GEN_15;
                                            end else begin
                                              if (6'h1a == _T_223) begin
                                                mem_26 <= _GEN_14;
                                              end else begin
                                                if (6'h1a == _T_218) begin
                                                  mem_26 <= _GEN_13;
                                                end else begin
                                                  if (6'h1a == _T_213) begin
                                                    mem_26 <= _GEN_12;
                                                  end else begin
                                                    if (6'h1a == _T_208) begin
                                                      mem_26 <= _GEN_11;
                                                    end else begin
                                                      if (6'h1a == _T_203) begin
                                                        mem_26 <= _GEN_10;
                                                      end else begin
                                                        if (6'h1a == _T_198) begin
                                                          mem_26 <= _GEN_9;
                                                        end else begin
                                                          if (6'h1a == _T_193) begin
                                                            mem_26 <= _GEN_8;
                                                          end else begin
                                                            if (6'h1a == _T_188) begin
                                                              mem_26 <= _GEN_7;
                                                            end else begin
                                                              if (6'h1a == _T_183) begin
                                                                mem_26 <= _GEN_6;
                                                              end else begin
                                                                if (6'h1a == _T_178) begin
                                                                  mem_26 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h1a == _T_173) begin
                                                                    mem_26 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h1a == _T_168) begin
                                                                      mem_26 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h1a == _T_163) begin
                                                                        mem_26 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h1a == _T_158) begin
                                                                          mem_26 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h1a == _T_153) begin
                                                                            mem_26 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h1a == _T_308) begin
            mem_26 <= _GEN_31;
          end else begin
            if (6'h1a == _T_303) begin
              mem_26 <= _GEN_30;
            end else begin
              if (6'h1a == _T_298) begin
                mem_26 <= _GEN_29;
              end else begin
                if (6'h1a == _T_293) begin
                  mem_26 <= _GEN_28;
                end else begin
                  if (6'h1a == _T_288) begin
                    mem_26 <= _GEN_27;
                  end else begin
                    if (6'h1a == _T_283) begin
                      mem_26 <= _GEN_26;
                    end else begin
                      if (6'h1a == _T_278) begin
                        mem_26 <= _GEN_25;
                      end else begin
                        if (6'h1a == _T_273) begin
                          mem_26 <= _GEN_24;
                        end else begin
                          if (6'h1a == _T_268) begin
                            mem_26 <= _GEN_23;
                          end else begin
                            if (6'h1a == _T_263) begin
                              mem_26 <= _GEN_22;
                            end else begin
                              if (6'h1a == _T_258) begin
                                mem_26 <= _GEN_21;
                              end else begin
                                if (6'h1a == _T_253) begin
                                  mem_26 <= _GEN_20;
                                end else begin
                                  if (6'h1a == _T_248) begin
                                    mem_26 <= _GEN_19;
                                  end else begin
                                    if (6'h1a == _T_243) begin
                                      mem_26 <= _GEN_18;
                                    end else begin
                                      if (6'h1a == _T_238) begin
                                        mem_26 <= _GEN_17;
                                      end else begin
                                        if (6'h1a == _T_233) begin
                                          mem_26 <= _GEN_16;
                                        end else begin
                                          if (6'h1a == _T_228) begin
                                            mem_26 <= _GEN_15;
                                          end else begin
                                            if (6'h1a == _T_223) begin
                                              mem_26 <= _GEN_14;
                                            end else begin
                                              if (6'h1a == _T_218) begin
                                                mem_26 <= _GEN_13;
                                              end else begin
                                                if (6'h1a == _T_213) begin
                                                  mem_26 <= _GEN_12;
                                                end else begin
                                                  if (6'h1a == _T_208) begin
                                                    mem_26 <= _GEN_11;
                                                  end else begin
                                                    if (6'h1a == _T_203) begin
                                                      mem_26 <= _GEN_10;
                                                    end else begin
                                                      if (6'h1a == _T_198) begin
                                                        mem_26 <= _GEN_9;
                                                      end else begin
                                                        if (6'h1a == _T_193) begin
                                                          mem_26 <= _GEN_8;
                                                        end else begin
                                                          if (6'h1a == _T_188) begin
                                                            mem_26 <= _GEN_7;
                                                          end else begin
                                                            if (6'h1a == _T_183) begin
                                                              mem_26 <= _GEN_6;
                                                            end else begin
                                                              if (6'h1a == _T_178) begin
                                                                mem_26 <= _GEN_5;
                                                              end else begin
                                                                if (6'h1a == _T_173) begin
                                                                  mem_26 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h1a == _T_168) begin
                                                                    mem_26 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h1a == _T_163) begin
                                                                      mem_26 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h1a == _T_158) begin
                                                                        mem_26 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h1a == _T_153) begin
                                                                          mem_26 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h1a == _T_308) begin
          mem_26 <= _GEN_31;
        end else begin
          if (6'h1a == _T_303) begin
            mem_26 <= _GEN_30;
          end else begin
            if (6'h1a == _T_298) begin
              mem_26 <= _GEN_29;
            end else begin
              if (6'h1a == _T_293) begin
                mem_26 <= _GEN_28;
              end else begin
                if (6'h1a == _T_288) begin
                  mem_26 <= _GEN_27;
                end else begin
                  if (6'h1a == _T_283) begin
                    mem_26 <= _GEN_26;
                  end else begin
                    if (6'h1a == _T_278) begin
                      mem_26 <= _GEN_25;
                    end else begin
                      if (6'h1a == _T_273) begin
                        mem_26 <= _GEN_24;
                      end else begin
                        if (6'h1a == _T_268) begin
                          mem_26 <= _GEN_23;
                        end else begin
                          if (6'h1a == _T_263) begin
                            mem_26 <= _GEN_22;
                          end else begin
                            if (6'h1a == _T_258) begin
                              mem_26 <= _GEN_21;
                            end else begin
                              if (6'h1a == _T_253) begin
                                mem_26 <= _GEN_20;
                              end else begin
                                if (6'h1a == _T_248) begin
                                  mem_26 <= _GEN_19;
                                end else begin
                                  if (6'h1a == _T_243) begin
                                    mem_26 <= _GEN_18;
                                  end else begin
                                    if (6'h1a == _T_238) begin
                                      mem_26 <= _GEN_17;
                                    end else begin
                                      if (6'h1a == _T_233) begin
                                        mem_26 <= _GEN_16;
                                      end else begin
                                        if (6'h1a == _T_228) begin
                                          mem_26 <= _GEN_15;
                                        end else begin
                                          if (6'h1a == _T_223) begin
                                            mem_26 <= _GEN_14;
                                          end else begin
                                            if (6'h1a == _T_218) begin
                                              mem_26 <= _GEN_13;
                                            end else begin
                                              if (6'h1a == _T_213) begin
                                                mem_26 <= _GEN_12;
                                              end else begin
                                                if (6'h1a == _T_208) begin
                                                  mem_26 <= _GEN_11;
                                                end else begin
                                                  if (6'h1a == _T_203) begin
                                                    mem_26 <= _GEN_10;
                                                  end else begin
                                                    if (6'h1a == _T_198) begin
                                                      mem_26 <= _GEN_9;
                                                    end else begin
                                                      if (6'h1a == _T_193) begin
                                                        mem_26 <= _GEN_8;
                                                      end else begin
                                                        if (6'h1a == _T_188) begin
                                                          mem_26 <= _GEN_7;
                                                        end else begin
                                                          if (6'h1a == _T_183) begin
                                                            mem_26 <= _GEN_6;
                                                          end else begin
                                                            if (6'h1a == _T_178) begin
                                                              mem_26 <= _GEN_5;
                                                            end else begin
                                                              if (6'h1a == _T_173) begin
                                                                mem_26 <= _GEN_4;
                                                              end else begin
                                                                if (6'h1a == _T_168) begin
                                                                  mem_26 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h1a == _T_163) begin
                                                                    mem_26 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h1a == _T_158) begin
                                                                      mem_26 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h1a == _T_153) begin
                                                                        mem_26 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h1b == wPos) begin
            mem_27 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h1b == _T_308) begin
                mem_27 <= _GEN_31;
              end else begin
                if (6'h1b == _T_303) begin
                  mem_27 <= _GEN_30;
                end else begin
                  if (6'h1b == _T_298) begin
                    mem_27 <= _GEN_29;
                  end else begin
                    if (6'h1b == _T_293) begin
                      mem_27 <= _GEN_28;
                    end else begin
                      if (6'h1b == _T_288) begin
                        mem_27 <= _GEN_27;
                      end else begin
                        if (6'h1b == _T_283) begin
                          mem_27 <= _GEN_26;
                        end else begin
                          if (6'h1b == _T_278) begin
                            mem_27 <= _GEN_25;
                          end else begin
                            if (6'h1b == _T_273) begin
                              mem_27 <= _GEN_24;
                            end else begin
                              if (6'h1b == _T_268) begin
                                mem_27 <= _GEN_23;
                              end else begin
                                if (6'h1b == _T_263) begin
                                  mem_27 <= _GEN_22;
                                end else begin
                                  if (6'h1b == _T_258) begin
                                    mem_27 <= _GEN_21;
                                  end else begin
                                    if (6'h1b == _T_253) begin
                                      mem_27 <= _GEN_20;
                                    end else begin
                                      if (6'h1b == _T_248) begin
                                        mem_27 <= _GEN_19;
                                      end else begin
                                        if (6'h1b == _T_243) begin
                                          mem_27 <= _GEN_18;
                                        end else begin
                                          if (6'h1b == _T_238) begin
                                            mem_27 <= _GEN_17;
                                          end else begin
                                            if (6'h1b == _T_233) begin
                                              mem_27 <= _GEN_16;
                                            end else begin
                                              if (6'h1b == _T_228) begin
                                                mem_27 <= _GEN_15;
                                              end else begin
                                                if (6'h1b == _T_223) begin
                                                  mem_27 <= _GEN_14;
                                                end else begin
                                                  if (6'h1b == _T_218) begin
                                                    mem_27 <= _GEN_13;
                                                  end else begin
                                                    if (6'h1b == _T_213) begin
                                                      mem_27 <= _GEN_12;
                                                    end else begin
                                                      if (6'h1b == _T_208) begin
                                                        mem_27 <= _GEN_11;
                                                      end else begin
                                                        if (6'h1b == _T_203) begin
                                                          mem_27 <= _GEN_10;
                                                        end else begin
                                                          if (6'h1b == _T_198) begin
                                                            mem_27 <= _GEN_9;
                                                          end else begin
                                                            if (6'h1b == _T_193) begin
                                                              mem_27 <= _GEN_8;
                                                            end else begin
                                                              if (6'h1b == _T_188) begin
                                                                mem_27 <= _GEN_7;
                                                              end else begin
                                                                if (6'h1b == _T_183) begin
                                                                  mem_27 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h1b == _T_178) begin
                                                                    mem_27 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h1b == _T_173) begin
                                                                      mem_27 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h1b == _T_168) begin
                                                                        mem_27 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h1b == _T_163) begin
                                                                          mem_27 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h1b == _T_158) begin
                                                                            mem_27 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h1b == _T_153) begin
                                                                              mem_27 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h1b == _T_308) begin
              mem_27 <= _GEN_31;
            end else begin
              if (6'h1b == _T_303) begin
                mem_27 <= _GEN_30;
              end else begin
                if (6'h1b == _T_298) begin
                  mem_27 <= _GEN_29;
                end else begin
                  if (6'h1b == _T_293) begin
                    mem_27 <= _GEN_28;
                  end else begin
                    if (6'h1b == _T_288) begin
                      mem_27 <= _GEN_27;
                    end else begin
                      if (6'h1b == _T_283) begin
                        mem_27 <= _GEN_26;
                      end else begin
                        if (6'h1b == _T_278) begin
                          mem_27 <= _GEN_25;
                        end else begin
                          if (6'h1b == _T_273) begin
                            mem_27 <= _GEN_24;
                          end else begin
                            if (6'h1b == _T_268) begin
                              mem_27 <= _GEN_23;
                            end else begin
                              if (6'h1b == _T_263) begin
                                mem_27 <= _GEN_22;
                              end else begin
                                if (6'h1b == _T_258) begin
                                  mem_27 <= _GEN_21;
                                end else begin
                                  if (6'h1b == _T_253) begin
                                    mem_27 <= _GEN_20;
                                  end else begin
                                    if (6'h1b == _T_248) begin
                                      mem_27 <= _GEN_19;
                                    end else begin
                                      if (6'h1b == _T_243) begin
                                        mem_27 <= _GEN_18;
                                      end else begin
                                        if (6'h1b == _T_238) begin
                                          mem_27 <= _GEN_17;
                                        end else begin
                                          if (6'h1b == _T_233) begin
                                            mem_27 <= _GEN_16;
                                          end else begin
                                            if (6'h1b == _T_228) begin
                                              mem_27 <= _GEN_15;
                                            end else begin
                                              if (6'h1b == _T_223) begin
                                                mem_27 <= _GEN_14;
                                              end else begin
                                                if (6'h1b == _T_218) begin
                                                  mem_27 <= _GEN_13;
                                                end else begin
                                                  if (6'h1b == _T_213) begin
                                                    mem_27 <= _GEN_12;
                                                  end else begin
                                                    if (6'h1b == _T_208) begin
                                                      mem_27 <= _GEN_11;
                                                    end else begin
                                                      if (6'h1b == _T_203) begin
                                                        mem_27 <= _GEN_10;
                                                      end else begin
                                                        if (6'h1b == _T_198) begin
                                                          mem_27 <= _GEN_9;
                                                        end else begin
                                                          if (6'h1b == _T_193) begin
                                                            mem_27 <= _GEN_8;
                                                          end else begin
                                                            if (6'h1b == _T_188) begin
                                                              mem_27 <= _GEN_7;
                                                            end else begin
                                                              if (6'h1b == _T_183) begin
                                                                mem_27 <= _GEN_6;
                                                              end else begin
                                                                if (6'h1b == _T_178) begin
                                                                  mem_27 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h1b == _T_173) begin
                                                                    mem_27 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h1b == _T_168) begin
                                                                      mem_27 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h1b == _T_163) begin
                                                                        mem_27 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h1b == _T_158) begin
                                                                          mem_27 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h1b == _T_153) begin
                                                                            mem_27 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h1b == _T_308) begin
            mem_27 <= _GEN_31;
          end else begin
            if (6'h1b == _T_303) begin
              mem_27 <= _GEN_30;
            end else begin
              if (6'h1b == _T_298) begin
                mem_27 <= _GEN_29;
              end else begin
                if (6'h1b == _T_293) begin
                  mem_27 <= _GEN_28;
                end else begin
                  if (6'h1b == _T_288) begin
                    mem_27 <= _GEN_27;
                  end else begin
                    if (6'h1b == _T_283) begin
                      mem_27 <= _GEN_26;
                    end else begin
                      if (6'h1b == _T_278) begin
                        mem_27 <= _GEN_25;
                      end else begin
                        if (6'h1b == _T_273) begin
                          mem_27 <= _GEN_24;
                        end else begin
                          if (6'h1b == _T_268) begin
                            mem_27 <= _GEN_23;
                          end else begin
                            if (6'h1b == _T_263) begin
                              mem_27 <= _GEN_22;
                            end else begin
                              if (6'h1b == _T_258) begin
                                mem_27 <= _GEN_21;
                              end else begin
                                if (6'h1b == _T_253) begin
                                  mem_27 <= _GEN_20;
                                end else begin
                                  if (6'h1b == _T_248) begin
                                    mem_27 <= _GEN_19;
                                  end else begin
                                    if (6'h1b == _T_243) begin
                                      mem_27 <= _GEN_18;
                                    end else begin
                                      if (6'h1b == _T_238) begin
                                        mem_27 <= _GEN_17;
                                      end else begin
                                        if (6'h1b == _T_233) begin
                                          mem_27 <= _GEN_16;
                                        end else begin
                                          if (6'h1b == _T_228) begin
                                            mem_27 <= _GEN_15;
                                          end else begin
                                            if (6'h1b == _T_223) begin
                                              mem_27 <= _GEN_14;
                                            end else begin
                                              if (6'h1b == _T_218) begin
                                                mem_27 <= _GEN_13;
                                              end else begin
                                                if (6'h1b == _T_213) begin
                                                  mem_27 <= _GEN_12;
                                                end else begin
                                                  if (6'h1b == _T_208) begin
                                                    mem_27 <= _GEN_11;
                                                  end else begin
                                                    if (6'h1b == _T_203) begin
                                                      mem_27 <= _GEN_10;
                                                    end else begin
                                                      if (6'h1b == _T_198) begin
                                                        mem_27 <= _GEN_9;
                                                      end else begin
                                                        if (6'h1b == _T_193) begin
                                                          mem_27 <= _GEN_8;
                                                        end else begin
                                                          if (6'h1b == _T_188) begin
                                                            mem_27 <= _GEN_7;
                                                          end else begin
                                                            if (6'h1b == _T_183) begin
                                                              mem_27 <= _GEN_6;
                                                            end else begin
                                                              if (6'h1b == _T_178) begin
                                                                mem_27 <= _GEN_5;
                                                              end else begin
                                                                if (6'h1b == _T_173) begin
                                                                  mem_27 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h1b == _T_168) begin
                                                                    mem_27 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h1b == _T_163) begin
                                                                      mem_27 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h1b == _T_158) begin
                                                                        mem_27 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h1b == _T_153) begin
                                                                          mem_27 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h1b == _T_308) begin
          mem_27 <= _GEN_31;
        end else begin
          if (6'h1b == _T_303) begin
            mem_27 <= _GEN_30;
          end else begin
            if (6'h1b == _T_298) begin
              mem_27 <= _GEN_29;
            end else begin
              if (6'h1b == _T_293) begin
                mem_27 <= _GEN_28;
              end else begin
                if (6'h1b == _T_288) begin
                  mem_27 <= _GEN_27;
                end else begin
                  if (6'h1b == _T_283) begin
                    mem_27 <= _GEN_26;
                  end else begin
                    if (6'h1b == _T_278) begin
                      mem_27 <= _GEN_25;
                    end else begin
                      if (6'h1b == _T_273) begin
                        mem_27 <= _GEN_24;
                      end else begin
                        if (6'h1b == _T_268) begin
                          mem_27 <= _GEN_23;
                        end else begin
                          if (6'h1b == _T_263) begin
                            mem_27 <= _GEN_22;
                          end else begin
                            if (6'h1b == _T_258) begin
                              mem_27 <= _GEN_21;
                            end else begin
                              if (6'h1b == _T_253) begin
                                mem_27 <= _GEN_20;
                              end else begin
                                if (6'h1b == _T_248) begin
                                  mem_27 <= _GEN_19;
                                end else begin
                                  if (6'h1b == _T_243) begin
                                    mem_27 <= _GEN_18;
                                  end else begin
                                    if (6'h1b == _T_238) begin
                                      mem_27 <= _GEN_17;
                                    end else begin
                                      if (6'h1b == _T_233) begin
                                        mem_27 <= _GEN_16;
                                      end else begin
                                        if (6'h1b == _T_228) begin
                                          mem_27 <= _GEN_15;
                                        end else begin
                                          if (6'h1b == _T_223) begin
                                            mem_27 <= _GEN_14;
                                          end else begin
                                            if (6'h1b == _T_218) begin
                                              mem_27 <= _GEN_13;
                                            end else begin
                                              if (6'h1b == _T_213) begin
                                                mem_27 <= _GEN_12;
                                              end else begin
                                                if (6'h1b == _T_208) begin
                                                  mem_27 <= _GEN_11;
                                                end else begin
                                                  if (6'h1b == _T_203) begin
                                                    mem_27 <= _GEN_10;
                                                  end else begin
                                                    if (6'h1b == _T_198) begin
                                                      mem_27 <= _GEN_9;
                                                    end else begin
                                                      if (6'h1b == _T_193) begin
                                                        mem_27 <= _GEN_8;
                                                      end else begin
                                                        if (6'h1b == _T_188) begin
                                                          mem_27 <= _GEN_7;
                                                        end else begin
                                                          if (6'h1b == _T_183) begin
                                                            mem_27 <= _GEN_6;
                                                          end else begin
                                                            if (6'h1b == _T_178) begin
                                                              mem_27 <= _GEN_5;
                                                            end else begin
                                                              if (6'h1b == _T_173) begin
                                                                mem_27 <= _GEN_4;
                                                              end else begin
                                                                if (6'h1b == _T_168) begin
                                                                  mem_27 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h1b == _T_163) begin
                                                                    mem_27 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h1b == _T_158) begin
                                                                      mem_27 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h1b == _T_153) begin
                                                                        mem_27 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h1c == wPos) begin
            mem_28 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h1c == _T_308) begin
                mem_28 <= _GEN_31;
              end else begin
                if (6'h1c == _T_303) begin
                  mem_28 <= _GEN_30;
                end else begin
                  if (6'h1c == _T_298) begin
                    mem_28 <= _GEN_29;
                  end else begin
                    if (6'h1c == _T_293) begin
                      mem_28 <= _GEN_28;
                    end else begin
                      if (6'h1c == _T_288) begin
                        mem_28 <= _GEN_27;
                      end else begin
                        if (6'h1c == _T_283) begin
                          mem_28 <= _GEN_26;
                        end else begin
                          if (6'h1c == _T_278) begin
                            mem_28 <= _GEN_25;
                          end else begin
                            if (6'h1c == _T_273) begin
                              mem_28 <= _GEN_24;
                            end else begin
                              if (6'h1c == _T_268) begin
                                mem_28 <= _GEN_23;
                              end else begin
                                if (6'h1c == _T_263) begin
                                  mem_28 <= _GEN_22;
                                end else begin
                                  if (6'h1c == _T_258) begin
                                    mem_28 <= _GEN_21;
                                  end else begin
                                    if (6'h1c == _T_253) begin
                                      mem_28 <= _GEN_20;
                                    end else begin
                                      if (6'h1c == _T_248) begin
                                        mem_28 <= _GEN_19;
                                      end else begin
                                        if (6'h1c == _T_243) begin
                                          mem_28 <= _GEN_18;
                                        end else begin
                                          if (6'h1c == _T_238) begin
                                            mem_28 <= _GEN_17;
                                          end else begin
                                            if (6'h1c == _T_233) begin
                                              mem_28 <= _GEN_16;
                                            end else begin
                                              if (6'h1c == _T_228) begin
                                                mem_28 <= _GEN_15;
                                              end else begin
                                                if (6'h1c == _T_223) begin
                                                  mem_28 <= _GEN_14;
                                                end else begin
                                                  if (6'h1c == _T_218) begin
                                                    mem_28 <= _GEN_13;
                                                  end else begin
                                                    if (6'h1c == _T_213) begin
                                                      mem_28 <= _GEN_12;
                                                    end else begin
                                                      if (6'h1c == _T_208) begin
                                                        mem_28 <= _GEN_11;
                                                      end else begin
                                                        if (6'h1c == _T_203) begin
                                                          mem_28 <= _GEN_10;
                                                        end else begin
                                                          if (6'h1c == _T_198) begin
                                                            mem_28 <= _GEN_9;
                                                          end else begin
                                                            if (6'h1c == _T_193) begin
                                                              mem_28 <= _GEN_8;
                                                            end else begin
                                                              if (6'h1c == _T_188) begin
                                                                mem_28 <= _GEN_7;
                                                              end else begin
                                                                if (6'h1c == _T_183) begin
                                                                  mem_28 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h1c == _T_178) begin
                                                                    mem_28 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h1c == _T_173) begin
                                                                      mem_28 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h1c == _T_168) begin
                                                                        mem_28 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h1c == _T_163) begin
                                                                          mem_28 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h1c == _T_158) begin
                                                                            mem_28 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h1c == _T_153) begin
                                                                              mem_28 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h1c == _T_308) begin
              mem_28 <= _GEN_31;
            end else begin
              if (6'h1c == _T_303) begin
                mem_28 <= _GEN_30;
              end else begin
                if (6'h1c == _T_298) begin
                  mem_28 <= _GEN_29;
                end else begin
                  if (6'h1c == _T_293) begin
                    mem_28 <= _GEN_28;
                  end else begin
                    if (6'h1c == _T_288) begin
                      mem_28 <= _GEN_27;
                    end else begin
                      if (6'h1c == _T_283) begin
                        mem_28 <= _GEN_26;
                      end else begin
                        if (6'h1c == _T_278) begin
                          mem_28 <= _GEN_25;
                        end else begin
                          if (6'h1c == _T_273) begin
                            mem_28 <= _GEN_24;
                          end else begin
                            if (6'h1c == _T_268) begin
                              mem_28 <= _GEN_23;
                            end else begin
                              if (6'h1c == _T_263) begin
                                mem_28 <= _GEN_22;
                              end else begin
                                if (6'h1c == _T_258) begin
                                  mem_28 <= _GEN_21;
                                end else begin
                                  if (6'h1c == _T_253) begin
                                    mem_28 <= _GEN_20;
                                  end else begin
                                    if (6'h1c == _T_248) begin
                                      mem_28 <= _GEN_19;
                                    end else begin
                                      if (6'h1c == _T_243) begin
                                        mem_28 <= _GEN_18;
                                      end else begin
                                        if (6'h1c == _T_238) begin
                                          mem_28 <= _GEN_17;
                                        end else begin
                                          if (6'h1c == _T_233) begin
                                            mem_28 <= _GEN_16;
                                          end else begin
                                            if (6'h1c == _T_228) begin
                                              mem_28 <= _GEN_15;
                                            end else begin
                                              if (6'h1c == _T_223) begin
                                                mem_28 <= _GEN_14;
                                              end else begin
                                                if (6'h1c == _T_218) begin
                                                  mem_28 <= _GEN_13;
                                                end else begin
                                                  if (6'h1c == _T_213) begin
                                                    mem_28 <= _GEN_12;
                                                  end else begin
                                                    if (6'h1c == _T_208) begin
                                                      mem_28 <= _GEN_11;
                                                    end else begin
                                                      if (6'h1c == _T_203) begin
                                                        mem_28 <= _GEN_10;
                                                      end else begin
                                                        if (6'h1c == _T_198) begin
                                                          mem_28 <= _GEN_9;
                                                        end else begin
                                                          if (6'h1c == _T_193) begin
                                                            mem_28 <= _GEN_8;
                                                          end else begin
                                                            if (6'h1c == _T_188) begin
                                                              mem_28 <= _GEN_7;
                                                            end else begin
                                                              if (6'h1c == _T_183) begin
                                                                mem_28 <= _GEN_6;
                                                              end else begin
                                                                if (6'h1c == _T_178) begin
                                                                  mem_28 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h1c == _T_173) begin
                                                                    mem_28 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h1c == _T_168) begin
                                                                      mem_28 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h1c == _T_163) begin
                                                                        mem_28 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h1c == _T_158) begin
                                                                          mem_28 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h1c == _T_153) begin
                                                                            mem_28 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h1c == _T_308) begin
            mem_28 <= _GEN_31;
          end else begin
            if (6'h1c == _T_303) begin
              mem_28 <= _GEN_30;
            end else begin
              if (6'h1c == _T_298) begin
                mem_28 <= _GEN_29;
              end else begin
                if (6'h1c == _T_293) begin
                  mem_28 <= _GEN_28;
                end else begin
                  if (6'h1c == _T_288) begin
                    mem_28 <= _GEN_27;
                  end else begin
                    if (6'h1c == _T_283) begin
                      mem_28 <= _GEN_26;
                    end else begin
                      if (6'h1c == _T_278) begin
                        mem_28 <= _GEN_25;
                      end else begin
                        if (6'h1c == _T_273) begin
                          mem_28 <= _GEN_24;
                        end else begin
                          if (6'h1c == _T_268) begin
                            mem_28 <= _GEN_23;
                          end else begin
                            if (6'h1c == _T_263) begin
                              mem_28 <= _GEN_22;
                            end else begin
                              if (6'h1c == _T_258) begin
                                mem_28 <= _GEN_21;
                              end else begin
                                if (6'h1c == _T_253) begin
                                  mem_28 <= _GEN_20;
                                end else begin
                                  if (6'h1c == _T_248) begin
                                    mem_28 <= _GEN_19;
                                  end else begin
                                    if (6'h1c == _T_243) begin
                                      mem_28 <= _GEN_18;
                                    end else begin
                                      if (6'h1c == _T_238) begin
                                        mem_28 <= _GEN_17;
                                      end else begin
                                        if (6'h1c == _T_233) begin
                                          mem_28 <= _GEN_16;
                                        end else begin
                                          if (6'h1c == _T_228) begin
                                            mem_28 <= _GEN_15;
                                          end else begin
                                            if (6'h1c == _T_223) begin
                                              mem_28 <= _GEN_14;
                                            end else begin
                                              if (6'h1c == _T_218) begin
                                                mem_28 <= _GEN_13;
                                              end else begin
                                                if (6'h1c == _T_213) begin
                                                  mem_28 <= _GEN_12;
                                                end else begin
                                                  if (6'h1c == _T_208) begin
                                                    mem_28 <= _GEN_11;
                                                  end else begin
                                                    if (6'h1c == _T_203) begin
                                                      mem_28 <= _GEN_10;
                                                    end else begin
                                                      if (6'h1c == _T_198) begin
                                                        mem_28 <= _GEN_9;
                                                      end else begin
                                                        if (6'h1c == _T_193) begin
                                                          mem_28 <= _GEN_8;
                                                        end else begin
                                                          if (6'h1c == _T_188) begin
                                                            mem_28 <= _GEN_7;
                                                          end else begin
                                                            if (6'h1c == _T_183) begin
                                                              mem_28 <= _GEN_6;
                                                            end else begin
                                                              if (6'h1c == _T_178) begin
                                                                mem_28 <= _GEN_5;
                                                              end else begin
                                                                if (6'h1c == _T_173) begin
                                                                  mem_28 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h1c == _T_168) begin
                                                                    mem_28 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h1c == _T_163) begin
                                                                      mem_28 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h1c == _T_158) begin
                                                                        mem_28 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h1c == _T_153) begin
                                                                          mem_28 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h1c == _T_308) begin
          mem_28 <= _GEN_31;
        end else begin
          if (6'h1c == _T_303) begin
            mem_28 <= _GEN_30;
          end else begin
            if (6'h1c == _T_298) begin
              mem_28 <= _GEN_29;
            end else begin
              if (6'h1c == _T_293) begin
                mem_28 <= _GEN_28;
              end else begin
                if (6'h1c == _T_288) begin
                  mem_28 <= _GEN_27;
                end else begin
                  if (6'h1c == _T_283) begin
                    mem_28 <= _GEN_26;
                  end else begin
                    if (6'h1c == _T_278) begin
                      mem_28 <= _GEN_25;
                    end else begin
                      if (6'h1c == _T_273) begin
                        mem_28 <= _GEN_24;
                      end else begin
                        if (6'h1c == _T_268) begin
                          mem_28 <= _GEN_23;
                        end else begin
                          if (6'h1c == _T_263) begin
                            mem_28 <= _GEN_22;
                          end else begin
                            if (6'h1c == _T_258) begin
                              mem_28 <= _GEN_21;
                            end else begin
                              if (6'h1c == _T_253) begin
                                mem_28 <= _GEN_20;
                              end else begin
                                if (6'h1c == _T_248) begin
                                  mem_28 <= _GEN_19;
                                end else begin
                                  if (6'h1c == _T_243) begin
                                    mem_28 <= _GEN_18;
                                  end else begin
                                    if (6'h1c == _T_238) begin
                                      mem_28 <= _GEN_17;
                                    end else begin
                                      if (6'h1c == _T_233) begin
                                        mem_28 <= _GEN_16;
                                      end else begin
                                        if (6'h1c == _T_228) begin
                                          mem_28 <= _GEN_15;
                                        end else begin
                                          if (6'h1c == _T_223) begin
                                            mem_28 <= _GEN_14;
                                          end else begin
                                            if (6'h1c == _T_218) begin
                                              mem_28 <= _GEN_13;
                                            end else begin
                                              if (6'h1c == _T_213) begin
                                                mem_28 <= _GEN_12;
                                              end else begin
                                                if (6'h1c == _T_208) begin
                                                  mem_28 <= _GEN_11;
                                                end else begin
                                                  if (6'h1c == _T_203) begin
                                                    mem_28 <= _GEN_10;
                                                  end else begin
                                                    if (6'h1c == _T_198) begin
                                                      mem_28 <= _GEN_9;
                                                    end else begin
                                                      if (6'h1c == _T_193) begin
                                                        mem_28 <= _GEN_8;
                                                      end else begin
                                                        if (6'h1c == _T_188) begin
                                                          mem_28 <= _GEN_7;
                                                        end else begin
                                                          if (6'h1c == _T_183) begin
                                                            mem_28 <= _GEN_6;
                                                          end else begin
                                                            if (6'h1c == _T_178) begin
                                                              mem_28 <= _GEN_5;
                                                            end else begin
                                                              if (6'h1c == _T_173) begin
                                                                mem_28 <= _GEN_4;
                                                              end else begin
                                                                if (6'h1c == _T_168) begin
                                                                  mem_28 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h1c == _T_163) begin
                                                                    mem_28 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h1c == _T_158) begin
                                                                      mem_28 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h1c == _T_153) begin
                                                                        mem_28 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h1d == wPos) begin
            mem_29 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h1d == _T_308) begin
                mem_29 <= _GEN_31;
              end else begin
                if (6'h1d == _T_303) begin
                  mem_29 <= _GEN_30;
                end else begin
                  if (6'h1d == _T_298) begin
                    mem_29 <= _GEN_29;
                  end else begin
                    if (6'h1d == _T_293) begin
                      mem_29 <= _GEN_28;
                    end else begin
                      if (6'h1d == _T_288) begin
                        mem_29 <= _GEN_27;
                      end else begin
                        if (6'h1d == _T_283) begin
                          mem_29 <= _GEN_26;
                        end else begin
                          if (6'h1d == _T_278) begin
                            mem_29 <= _GEN_25;
                          end else begin
                            if (6'h1d == _T_273) begin
                              mem_29 <= _GEN_24;
                            end else begin
                              if (6'h1d == _T_268) begin
                                mem_29 <= _GEN_23;
                              end else begin
                                if (6'h1d == _T_263) begin
                                  mem_29 <= _GEN_22;
                                end else begin
                                  if (6'h1d == _T_258) begin
                                    mem_29 <= _GEN_21;
                                  end else begin
                                    if (6'h1d == _T_253) begin
                                      mem_29 <= _GEN_20;
                                    end else begin
                                      if (6'h1d == _T_248) begin
                                        mem_29 <= _GEN_19;
                                      end else begin
                                        if (6'h1d == _T_243) begin
                                          mem_29 <= _GEN_18;
                                        end else begin
                                          if (6'h1d == _T_238) begin
                                            mem_29 <= _GEN_17;
                                          end else begin
                                            if (6'h1d == _T_233) begin
                                              mem_29 <= _GEN_16;
                                            end else begin
                                              if (6'h1d == _T_228) begin
                                                mem_29 <= _GEN_15;
                                              end else begin
                                                if (6'h1d == _T_223) begin
                                                  mem_29 <= _GEN_14;
                                                end else begin
                                                  if (6'h1d == _T_218) begin
                                                    mem_29 <= _GEN_13;
                                                  end else begin
                                                    if (6'h1d == _T_213) begin
                                                      mem_29 <= _GEN_12;
                                                    end else begin
                                                      if (6'h1d == _T_208) begin
                                                        mem_29 <= _GEN_11;
                                                      end else begin
                                                        if (6'h1d == _T_203) begin
                                                          mem_29 <= _GEN_10;
                                                        end else begin
                                                          if (6'h1d == _T_198) begin
                                                            mem_29 <= _GEN_9;
                                                          end else begin
                                                            if (6'h1d == _T_193) begin
                                                              mem_29 <= _GEN_8;
                                                            end else begin
                                                              if (6'h1d == _T_188) begin
                                                                mem_29 <= _GEN_7;
                                                              end else begin
                                                                if (6'h1d == _T_183) begin
                                                                  mem_29 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h1d == _T_178) begin
                                                                    mem_29 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h1d == _T_173) begin
                                                                      mem_29 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h1d == _T_168) begin
                                                                        mem_29 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h1d == _T_163) begin
                                                                          mem_29 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h1d == _T_158) begin
                                                                            mem_29 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h1d == _T_153) begin
                                                                              mem_29 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h1d == _T_308) begin
              mem_29 <= _GEN_31;
            end else begin
              if (6'h1d == _T_303) begin
                mem_29 <= _GEN_30;
              end else begin
                if (6'h1d == _T_298) begin
                  mem_29 <= _GEN_29;
                end else begin
                  if (6'h1d == _T_293) begin
                    mem_29 <= _GEN_28;
                  end else begin
                    if (6'h1d == _T_288) begin
                      mem_29 <= _GEN_27;
                    end else begin
                      if (6'h1d == _T_283) begin
                        mem_29 <= _GEN_26;
                      end else begin
                        if (6'h1d == _T_278) begin
                          mem_29 <= _GEN_25;
                        end else begin
                          if (6'h1d == _T_273) begin
                            mem_29 <= _GEN_24;
                          end else begin
                            if (6'h1d == _T_268) begin
                              mem_29 <= _GEN_23;
                            end else begin
                              if (6'h1d == _T_263) begin
                                mem_29 <= _GEN_22;
                              end else begin
                                if (6'h1d == _T_258) begin
                                  mem_29 <= _GEN_21;
                                end else begin
                                  if (6'h1d == _T_253) begin
                                    mem_29 <= _GEN_20;
                                  end else begin
                                    if (6'h1d == _T_248) begin
                                      mem_29 <= _GEN_19;
                                    end else begin
                                      if (6'h1d == _T_243) begin
                                        mem_29 <= _GEN_18;
                                      end else begin
                                        if (6'h1d == _T_238) begin
                                          mem_29 <= _GEN_17;
                                        end else begin
                                          if (6'h1d == _T_233) begin
                                            mem_29 <= _GEN_16;
                                          end else begin
                                            if (6'h1d == _T_228) begin
                                              mem_29 <= _GEN_15;
                                            end else begin
                                              if (6'h1d == _T_223) begin
                                                mem_29 <= _GEN_14;
                                              end else begin
                                                if (6'h1d == _T_218) begin
                                                  mem_29 <= _GEN_13;
                                                end else begin
                                                  if (6'h1d == _T_213) begin
                                                    mem_29 <= _GEN_12;
                                                  end else begin
                                                    if (6'h1d == _T_208) begin
                                                      mem_29 <= _GEN_11;
                                                    end else begin
                                                      if (6'h1d == _T_203) begin
                                                        mem_29 <= _GEN_10;
                                                      end else begin
                                                        if (6'h1d == _T_198) begin
                                                          mem_29 <= _GEN_9;
                                                        end else begin
                                                          if (6'h1d == _T_193) begin
                                                            mem_29 <= _GEN_8;
                                                          end else begin
                                                            if (6'h1d == _T_188) begin
                                                              mem_29 <= _GEN_7;
                                                            end else begin
                                                              if (6'h1d == _T_183) begin
                                                                mem_29 <= _GEN_6;
                                                              end else begin
                                                                if (6'h1d == _T_178) begin
                                                                  mem_29 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h1d == _T_173) begin
                                                                    mem_29 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h1d == _T_168) begin
                                                                      mem_29 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h1d == _T_163) begin
                                                                        mem_29 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h1d == _T_158) begin
                                                                          mem_29 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h1d == _T_153) begin
                                                                            mem_29 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h1d == _T_308) begin
            mem_29 <= _GEN_31;
          end else begin
            if (6'h1d == _T_303) begin
              mem_29 <= _GEN_30;
            end else begin
              if (6'h1d == _T_298) begin
                mem_29 <= _GEN_29;
              end else begin
                if (6'h1d == _T_293) begin
                  mem_29 <= _GEN_28;
                end else begin
                  if (6'h1d == _T_288) begin
                    mem_29 <= _GEN_27;
                  end else begin
                    if (6'h1d == _T_283) begin
                      mem_29 <= _GEN_26;
                    end else begin
                      if (6'h1d == _T_278) begin
                        mem_29 <= _GEN_25;
                      end else begin
                        if (6'h1d == _T_273) begin
                          mem_29 <= _GEN_24;
                        end else begin
                          if (6'h1d == _T_268) begin
                            mem_29 <= _GEN_23;
                          end else begin
                            if (6'h1d == _T_263) begin
                              mem_29 <= _GEN_22;
                            end else begin
                              if (6'h1d == _T_258) begin
                                mem_29 <= _GEN_21;
                              end else begin
                                if (6'h1d == _T_253) begin
                                  mem_29 <= _GEN_20;
                                end else begin
                                  if (6'h1d == _T_248) begin
                                    mem_29 <= _GEN_19;
                                  end else begin
                                    if (6'h1d == _T_243) begin
                                      mem_29 <= _GEN_18;
                                    end else begin
                                      if (6'h1d == _T_238) begin
                                        mem_29 <= _GEN_17;
                                      end else begin
                                        if (6'h1d == _T_233) begin
                                          mem_29 <= _GEN_16;
                                        end else begin
                                          if (6'h1d == _T_228) begin
                                            mem_29 <= _GEN_15;
                                          end else begin
                                            if (6'h1d == _T_223) begin
                                              mem_29 <= _GEN_14;
                                            end else begin
                                              if (6'h1d == _T_218) begin
                                                mem_29 <= _GEN_13;
                                              end else begin
                                                if (6'h1d == _T_213) begin
                                                  mem_29 <= _GEN_12;
                                                end else begin
                                                  if (6'h1d == _T_208) begin
                                                    mem_29 <= _GEN_11;
                                                  end else begin
                                                    if (6'h1d == _T_203) begin
                                                      mem_29 <= _GEN_10;
                                                    end else begin
                                                      if (6'h1d == _T_198) begin
                                                        mem_29 <= _GEN_9;
                                                      end else begin
                                                        if (6'h1d == _T_193) begin
                                                          mem_29 <= _GEN_8;
                                                        end else begin
                                                          if (6'h1d == _T_188) begin
                                                            mem_29 <= _GEN_7;
                                                          end else begin
                                                            if (6'h1d == _T_183) begin
                                                              mem_29 <= _GEN_6;
                                                            end else begin
                                                              if (6'h1d == _T_178) begin
                                                                mem_29 <= _GEN_5;
                                                              end else begin
                                                                if (6'h1d == _T_173) begin
                                                                  mem_29 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h1d == _T_168) begin
                                                                    mem_29 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h1d == _T_163) begin
                                                                      mem_29 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h1d == _T_158) begin
                                                                        mem_29 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h1d == _T_153) begin
                                                                          mem_29 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h1d == _T_308) begin
          mem_29 <= _GEN_31;
        end else begin
          if (6'h1d == _T_303) begin
            mem_29 <= _GEN_30;
          end else begin
            if (6'h1d == _T_298) begin
              mem_29 <= _GEN_29;
            end else begin
              if (6'h1d == _T_293) begin
                mem_29 <= _GEN_28;
              end else begin
                if (6'h1d == _T_288) begin
                  mem_29 <= _GEN_27;
                end else begin
                  if (6'h1d == _T_283) begin
                    mem_29 <= _GEN_26;
                  end else begin
                    if (6'h1d == _T_278) begin
                      mem_29 <= _GEN_25;
                    end else begin
                      if (6'h1d == _T_273) begin
                        mem_29 <= _GEN_24;
                      end else begin
                        if (6'h1d == _T_268) begin
                          mem_29 <= _GEN_23;
                        end else begin
                          if (6'h1d == _T_263) begin
                            mem_29 <= _GEN_22;
                          end else begin
                            if (6'h1d == _T_258) begin
                              mem_29 <= _GEN_21;
                            end else begin
                              if (6'h1d == _T_253) begin
                                mem_29 <= _GEN_20;
                              end else begin
                                if (6'h1d == _T_248) begin
                                  mem_29 <= _GEN_19;
                                end else begin
                                  if (6'h1d == _T_243) begin
                                    mem_29 <= _GEN_18;
                                  end else begin
                                    if (6'h1d == _T_238) begin
                                      mem_29 <= _GEN_17;
                                    end else begin
                                      if (6'h1d == _T_233) begin
                                        mem_29 <= _GEN_16;
                                      end else begin
                                        if (6'h1d == _T_228) begin
                                          mem_29 <= _GEN_15;
                                        end else begin
                                          if (6'h1d == _T_223) begin
                                            mem_29 <= _GEN_14;
                                          end else begin
                                            if (6'h1d == _T_218) begin
                                              mem_29 <= _GEN_13;
                                            end else begin
                                              if (6'h1d == _T_213) begin
                                                mem_29 <= _GEN_12;
                                              end else begin
                                                if (6'h1d == _T_208) begin
                                                  mem_29 <= _GEN_11;
                                                end else begin
                                                  if (6'h1d == _T_203) begin
                                                    mem_29 <= _GEN_10;
                                                  end else begin
                                                    if (6'h1d == _T_198) begin
                                                      mem_29 <= _GEN_9;
                                                    end else begin
                                                      if (6'h1d == _T_193) begin
                                                        mem_29 <= _GEN_8;
                                                      end else begin
                                                        if (6'h1d == _T_188) begin
                                                          mem_29 <= _GEN_7;
                                                        end else begin
                                                          if (6'h1d == _T_183) begin
                                                            mem_29 <= _GEN_6;
                                                          end else begin
                                                            if (6'h1d == _T_178) begin
                                                              mem_29 <= _GEN_5;
                                                            end else begin
                                                              if (6'h1d == _T_173) begin
                                                                mem_29 <= _GEN_4;
                                                              end else begin
                                                                if (6'h1d == _T_168) begin
                                                                  mem_29 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h1d == _T_163) begin
                                                                    mem_29 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h1d == _T_158) begin
                                                                      mem_29 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h1d == _T_153) begin
                                                                        mem_29 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h1e == wPos) begin
            mem_30 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h1e == _T_308) begin
                mem_30 <= _GEN_31;
              end else begin
                if (6'h1e == _T_303) begin
                  mem_30 <= _GEN_30;
                end else begin
                  if (6'h1e == _T_298) begin
                    mem_30 <= _GEN_29;
                  end else begin
                    if (6'h1e == _T_293) begin
                      mem_30 <= _GEN_28;
                    end else begin
                      if (6'h1e == _T_288) begin
                        mem_30 <= _GEN_27;
                      end else begin
                        if (6'h1e == _T_283) begin
                          mem_30 <= _GEN_26;
                        end else begin
                          if (6'h1e == _T_278) begin
                            mem_30 <= _GEN_25;
                          end else begin
                            if (6'h1e == _T_273) begin
                              mem_30 <= _GEN_24;
                            end else begin
                              if (6'h1e == _T_268) begin
                                mem_30 <= _GEN_23;
                              end else begin
                                if (6'h1e == _T_263) begin
                                  mem_30 <= _GEN_22;
                                end else begin
                                  if (6'h1e == _T_258) begin
                                    mem_30 <= _GEN_21;
                                  end else begin
                                    if (6'h1e == _T_253) begin
                                      mem_30 <= _GEN_20;
                                    end else begin
                                      if (6'h1e == _T_248) begin
                                        mem_30 <= _GEN_19;
                                      end else begin
                                        if (6'h1e == _T_243) begin
                                          mem_30 <= _GEN_18;
                                        end else begin
                                          if (6'h1e == _T_238) begin
                                            mem_30 <= _GEN_17;
                                          end else begin
                                            if (6'h1e == _T_233) begin
                                              mem_30 <= _GEN_16;
                                            end else begin
                                              if (6'h1e == _T_228) begin
                                                mem_30 <= _GEN_15;
                                              end else begin
                                                if (6'h1e == _T_223) begin
                                                  mem_30 <= _GEN_14;
                                                end else begin
                                                  if (6'h1e == _T_218) begin
                                                    mem_30 <= _GEN_13;
                                                  end else begin
                                                    if (6'h1e == _T_213) begin
                                                      mem_30 <= _GEN_12;
                                                    end else begin
                                                      if (6'h1e == _T_208) begin
                                                        mem_30 <= _GEN_11;
                                                      end else begin
                                                        if (6'h1e == _T_203) begin
                                                          mem_30 <= _GEN_10;
                                                        end else begin
                                                          if (6'h1e == _T_198) begin
                                                            mem_30 <= _GEN_9;
                                                          end else begin
                                                            if (6'h1e == _T_193) begin
                                                              mem_30 <= _GEN_8;
                                                            end else begin
                                                              if (6'h1e == _T_188) begin
                                                                mem_30 <= _GEN_7;
                                                              end else begin
                                                                if (6'h1e == _T_183) begin
                                                                  mem_30 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h1e == _T_178) begin
                                                                    mem_30 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h1e == _T_173) begin
                                                                      mem_30 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h1e == _T_168) begin
                                                                        mem_30 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h1e == _T_163) begin
                                                                          mem_30 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h1e == _T_158) begin
                                                                            mem_30 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h1e == _T_153) begin
                                                                              mem_30 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h1e == _T_308) begin
              mem_30 <= _GEN_31;
            end else begin
              if (6'h1e == _T_303) begin
                mem_30 <= _GEN_30;
              end else begin
                if (6'h1e == _T_298) begin
                  mem_30 <= _GEN_29;
                end else begin
                  if (6'h1e == _T_293) begin
                    mem_30 <= _GEN_28;
                  end else begin
                    if (6'h1e == _T_288) begin
                      mem_30 <= _GEN_27;
                    end else begin
                      if (6'h1e == _T_283) begin
                        mem_30 <= _GEN_26;
                      end else begin
                        if (6'h1e == _T_278) begin
                          mem_30 <= _GEN_25;
                        end else begin
                          if (6'h1e == _T_273) begin
                            mem_30 <= _GEN_24;
                          end else begin
                            if (6'h1e == _T_268) begin
                              mem_30 <= _GEN_23;
                            end else begin
                              if (6'h1e == _T_263) begin
                                mem_30 <= _GEN_22;
                              end else begin
                                if (6'h1e == _T_258) begin
                                  mem_30 <= _GEN_21;
                                end else begin
                                  if (6'h1e == _T_253) begin
                                    mem_30 <= _GEN_20;
                                  end else begin
                                    if (6'h1e == _T_248) begin
                                      mem_30 <= _GEN_19;
                                    end else begin
                                      if (6'h1e == _T_243) begin
                                        mem_30 <= _GEN_18;
                                      end else begin
                                        if (6'h1e == _T_238) begin
                                          mem_30 <= _GEN_17;
                                        end else begin
                                          if (6'h1e == _T_233) begin
                                            mem_30 <= _GEN_16;
                                          end else begin
                                            if (6'h1e == _T_228) begin
                                              mem_30 <= _GEN_15;
                                            end else begin
                                              if (6'h1e == _T_223) begin
                                                mem_30 <= _GEN_14;
                                              end else begin
                                                if (6'h1e == _T_218) begin
                                                  mem_30 <= _GEN_13;
                                                end else begin
                                                  if (6'h1e == _T_213) begin
                                                    mem_30 <= _GEN_12;
                                                  end else begin
                                                    if (6'h1e == _T_208) begin
                                                      mem_30 <= _GEN_11;
                                                    end else begin
                                                      if (6'h1e == _T_203) begin
                                                        mem_30 <= _GEN_10;
                                                      end else begin
                                                        if (6'h1e == _T_198) begin
                                                          mem_30 <= _GEN_9;
                                                        end else begin
                                                          if (6'h1e == _T_193) begin
                                                            mem_30 <= _GEN_8;
                                                          end else begin
                                                            if (6'h1e == _T_188) begin
                                                              mem_30 <= _GEN_7;
                                                            end else begin
                                                              if (6'h1e == _T_183) begin
                                                                mem_30 <= _GEN_6;
                                                              end else begin
                                                                if (6'h1e == _T_178) begin
                                                                  mem_30 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h1e == _T_173) begin
                                                                    mem_30 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h1e == _T_168) begin
                                                                      mem_30 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h1e == _T_163) begin
                                                                        mem_30 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h1e == _T_158) begin
                                                                          mem_30 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h1e == _T_153) begin
                                                                            mem_30 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h1e == _T_308) begin
            mem_30 <= _GEN_31;
          end else begin
            if (6'h1e == _T_303) begin
              mem_30 <= _GEN_30;
            end else begin
              if (6'h1e == _T_298) begin
                mem_30 <= _GEN_29;
              end else begin
                if (6'h1e == _T_293) begin
                  mem_30 <= _GEN_28;
                end else begin
                  if (6'h1e == _T_288) begin
                    mem_30 <= _GEN_27;
                  end else begin
                    if (6'h1e == _T_283) begin
                      mem_30 <= _GEN_26;
                    end else begin
                      if (6'h1e == _T_278) begin
                        mem_30 <= _GEN_25;
                      end else begin
                        if (6'h1e == _T_273) begin
                          mem_30 <= _GEN_24;
                        end else begin
                          if (6'h1e == _T_268) begin
                            mem_30 <= _GEN_23;
                          end else begin
                            if (6'h1e == _T_263) begin
                              mem_30 <= _GEN_22;
                            end else begin
                              if (6'h1e == _T_258) begin
                                mem_30 <= _GEN_21;
                              end else begin
                                if (6'h1e == _T_253) begin
                                  mem_30 <= _GEN_20;
                                end else begin
                                  if (6'h1e == _T_248) begin
                                    mem_30 <= _GEN_19;
                                  end else begin
                                    if (6'h1e == _T_243) begin
                                      mem_30 <= _GEN_18;
                                    end else begin
                                      if (6'h1e == _T_238) begin
                                        mem_30 <= _GEN_17;
                                      end else begin
                                        if (6'h1e == _T_233) begin
                                          mem_30 <= _GEN_16;
                                        end else begin
                                          if (6'h1e == _T_228) begin
                                            mem_30 <= _GEN_15;
                                          end else begin
                                            if (6'h1e == _T_223) begin
                                              mem_30 <= _GEN_14;
                                            end else begin
                                              if (6'h1e == _T_218) begin
                                                mem_30 <= _GEN_13;
                                              end else begin
                                                if (6'h1e == _T_213) begin
                                                  mem_30 <= _GEN_12;
                                                end else begin
                                                  if (6'h1e == _T_208) begin
                                                    mem_30 <= _GEN_11;
                                                  end else begin
                                                    if (6'h1e == _T_203) begin
                                                      mem_30 <= _GEN_10;
                                                    end else begin
                                                      if (6'h1e == _T_198) begin
                                                        mem_30 <= _GEN_9;
                                                      end else begin
                                                        if (6'h1e == _T_193) begin
                                                          mem_30 <= _GEN_8;
                                                        end else begin
                                                          if (6'h1e == _T_188) begin
                                                            mem_30 <= _GEN_7;
                                                          end else begin
                                                            if (6'h1e == _T_183) begin
                                                              mem_30 <= _GEN_6;
                                                            end else begin
                                                              if (6'h1e == _T_178) begin
                                                                mem_30 <= _GEN_5;
                                                              end else begin
                                                                if (6'h1e == _T_173) begin
                                                                  mem_30 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h1e == _T_168) begin
                                                                    mem_30 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h1e == _T_163) begin
                                                                      mem_30 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h1e == _T_158) begin
                                                                        mem_30 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h1e == _T_153) begin
                                                                          mem_30 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h1e == _T_308) begin
          mem_30 <= _GEN_31;
        end else begin
          if (6'h1e == _T_303) begin
            mem_30 <= _GEN_30;
          end else begin
            if (6'h1e == _T_298) begin
              mem_30 <= _GEN_29;
            end else begin
              if (6'h1e == _T_293) begin
                mem_30 <= _GEN_28;
              end else begin
                if (6'h1e == _T_288) begin
                  mem_30 <= _GEN_27;
                end else begin
                  if (6'h1e == _T_283) begin
                    mem_30 <= _GEN_26;
                  end else begin
                    if (6'h1e == _T_278) begin
                      mem_30 <= _GEN_25;
                    end else begin
                      if (6'h1e == _T_273) begin
                        mem_30 <= _GEN_24;
                      end else begin
                        if (6'h1e == _T_268) begin
                          mem_30 <= _GEN_23;
                        end else begin
                          if (6'h1e == _T_263) begin
                            mem_30 <= _GEN_22;
                          end else begin
                            if (6'h1e == _T_258) begin
                              mem_30 <= _GEN_21;
                            end else begin
                              if (6'h1e == _T_253) begin
                                mem_30 <= _GEN_20;
                              end else begin
                                if (6'h1e == _T_248) begin
                                  mem_30 <= _GEN_19;
                                end else begin
                                  if (6'h1e == _T_243) begin
                                    mem_30 <= _GEN_18;
                                  end else begin
                                    if (6'h1e == _T_238) begin
                                      mem_30 <= _GEN_17;
                                    end else begin
                                      if (6'h1e == _T_233) begin
                                        mem_30 <= _GEN_16;
                                      end else begin
                                        if (6'h1e == _T_228) begin
                                          mem_30 <= _GEN_15;
                                        end else begin
                                          if (6'h1e == _T_223) begin
                                            mem_30 <= _GEN_14;
                                          end else begin
                                            if (6'h1e == _T_218) begin
                                              mem_30 <= _GEN_13;
                                            end else begin
                                              if (6'h1e == _T_213) begin
                                                mem_30 <= _GEN_12;
                                              end else begin
                                                if (6'h1e == _T_208) begin
                                                  mem_30 <= _GEN_11;
                                                end else begin
                                                  if (6'h1e == _T_203) begin
                                                    mem_30 <= _GEN_10;
                                                  end else begin
                                                    if (6'h1e == _T_198) begin
                                                      mem_30 <= _GEN_9;
                                                    end else begin
                                                      if (6'h1e == _T_193) begin
                                                        mem_30 <= _GEN_8;
                                                      end else begin
                                                        if (6'h1e == _T_188) begin
                                                          mem_30 <= _GEN_7;
                                                        end else begin
                                                          if (6'h1e == _T_183) begin
                                                            mem_30 <= _GEN_6;
                                                          end else begin
                                                            if (6'h1e == _T_178) begin
                                                              mem_30 <= _GEN_5;
                                                            end else begin
                                                              if (6'h1e == _T_173) begin
                                                                mem_30 <= _GEN_4;
                                                              end else begin
                                                                if (6'h1e == _T_168) begin
                                                                  mem_30 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h1e == _T_163) begin
                                                                    mem_30 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h1e == _T_158) begin
                                                                      mem_30 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h1e == _T_153) begin
                                                                        mem_30 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h1f == wPos) begin
            mem_31 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h1f == _T_308) begin
                mem_31 <= _GEN_31;
              end else begin
                if (6'h1f == _T_303) begin
                  mem_31 <= _GEN_30;
                end else begin
                  if (6'h1f == _T_298) begin
                    mem_31 <= _GEN_29;
                  end else begin
                    if (6'h1f == _T_293) begin
                      mem_31 <= _GEN_28;
                    end else begin
                      if (6'h1f == _T_288) begin
                        mem_31 <= _GEN_27;
                      end else begin
                        if (6'h1f == _T_283) begin
                          mem_31 <= _GEN_26;
                        end else begin
                          if (6'h1f == _T_278) begin
                            mem_31 <= _GEN_25;
                          end else begin
                            if (6'h1f == _T_273) begin
                              mem_31 <= _GEN_24;
                            end else begin
                              if (6'h1f == _T_268) begin
                                mem_31 <= _GEN_23;
                              end else begin
                                if (6'h1f == _T_263) begin
                                  mem_31 <= _GEN_22;
                                end else begin
                                  if (6'h1f == _T_258) begin
                                    mem_31 <= _GEN_21;
                                  end else begin
                                    if (6'h1f == _T_253) begin
                                      mem_31 <= _GEN_20;
                                    end else begin
                                      if (6'h1f == _T_248) begin
                                        mem_31 <= _GEN_19;
                                      end else begin
                                        if (6'h1f == _T_243) begin
                                          mem_31 <= _GEN_18;
                                        end else begin
                                          if (6'h1f == _T_238) begin
                                            mem_31 <= _GEN_17;
                                          end else begin
                                            if (6'h1f == _T_233) begin
                                              mem_31 <= _GEN_16;
                                            end else begin
                                              if (6'h1f == _T_228) begin
                                                mem_31 <= _GEN_15;
                                              end else begin
                                                if (6'h1f == _T_223) begin
                                                  mem_31 <= _GEN_14;
                                                end else begin
                                                  if (6'h1f == _T_218) begin
                                                    mem_31 <= _GEN_13;
                                                  end else begin
                                                    if (6'h1f == _T_213) begin
                                                      mem_31 <= _GEN_12;
                                                    end else begin
                                                      if (6'h1f == _T_208) begin
                                                        mem_31 <= _GEN_11;
                                                      end else begin
                                                        if (6'h1f == _T_203) begin
                                                          mem_31 <= _GEN_10;
                                                        end else begin
                                                          if (6'h1f == _T_198) begin
                                                            mem_31 <= _GEN_9;
                                                          end else begin
                                                            if (6'h1f == _T_193) begin
                                                              mem_31 <= _GEN_8;
                                                            end else begin
                                                              if (6'h1f == _T_188) begin
                                                                mem_31 <= _GEN_7;
                                                              end else begin
                                                                if (6'h1f == _T_183) begin
                                                                  mem_31 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h1f == _T_178) begin
                                                                    mem_31 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h1f == _T_173) begin
                                                                      mem_31 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h1f == _T_168) begin
                                                                        mem_31 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h1f == _T_163) begin
                                                                          mem_31 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h1f == _T_158) begin
                                                                            mem_31 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h1f == _T_153) begin
                                                                              mem_31 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h1f == _T_308) begin
              mem_31 <= _GEN_31;
            end else begin
              if (6'h1f == _T_303) begin
                mem_31 <= _GEN_30;
              end else begin
                if (6'h1f == _T_298) begin
                  mem_31 <= _GEN_29;
                end else begin
                  if (6'h1f == _T_293) begin
                    mem_31 <= _GEN_28;
                  end else begin
                    if (6'h1f == _T_288) begin
                      mem_31 <= _GEN_27;
                    end else begin
                      if (6'h1f == _T_283) begin
                        mem_31 <= _GEN_26;
                      end else begin
                        if (6'h1f == _T_278) begin
                          mem_31 <= _GEN_25;
                        end else begin
                          if (6'h1f == _T_273) begin
                            mem_31 <= _GEN_24;
                          end else begin
                            if (6'h1f == _T_268) begin
                              mem_31 <= _GEN_23;
                            end else begin
                              if (6'h1f == _T_263) begin
                                mem_31 <= _GEN_22;
                              end else begin
                                if (6'h1f == _T_258) begin
                                  mem_31 <= _GEN_21;
                                end else begin
                                  if (6'h1f == _T_253) begin
                                    mem_31 <= _GEN_20;
                                  end else begin
                                    if (6'h1f == _T_248) begin
                                      mem_31 <= _GEN_19;
                                    end else begin
                                      if (6'h1f == _T_243) begin
                                        mem_31 <= _GEN_18;
                                      end else begin
                                        if (6'h1f == _T_238) begin
                                          mem_31 <= _GEN_17;
                                        end else begin
                                          if (6'h1f == _T_233) begin
                                            mem_31 <= _GEN_16;
                                          end else begin
                                            if (6'h1f == _T_228) begin
                                              mem_31 <= _GEN_15;
                                            end else begin
                                              if (6'h1f == _T_223) begin
                                                mem_31 <= _GEN_14;
                                              end else begin
                                                if (6'h1f == _T_218) begin
                                                  mem_31 <= _GEN_13;
                                                end else begin
                                                  if (6'h1f == _T_213) begin
                                                    mem_31 <= _GEN_12;
                                                  end else begin
                                                    if (6'h1f == _T_208) begin
                                                      mem_31 <= _GEN_11;
                                                    end else begin
                                                      if (6'h1f == _T_203) begin
                                                        mem_31 <= _GEN_10;
                                                      end else begin
                                                        if (6'h1f == _T_198) begin
                                                          mem_31 <= _GEN_9;
                                                        end else begin
                                                          if (6'h1f == _T_193) begin
                                                            mem_31 <= _GEN_8;
                                                          end else begin
                                                            if (6'h1f == _T_188) begin
                                                              mem_31 <= _GEN_7;
                                                            end else begin
                                                              if (6'h1f == _T_183) begin
                                                                mem_31 <= _GEN_6;
                                                              end else begin
                                                                if (6'h1f == _T_178) begin
                                                                  mem_31 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h1f == _T_173) begin
                                                                    mem_31 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h1f == _T_168) begin
                                                                      mem_31 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h1f == _T_163) begin
                                                                        mem_31 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h1f == _T_158) begin
                                                                          mem_31 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h1f == _T_153) begin
                                                                            mem_31 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h1f == _T_308) begin
            mem_31 <= _GEN_31;
          end else begin
            if (6'h1f == _T_303) begin
              mem_31 <= _GEN_30;
            end else begin
              if (6'h1f == _T_298) begin
                mem_31 <= _GEN_29;
              end else begin
                if (6'h1f == _T_293) begin
                  mem_31 <= _GEN_28;
                end else begin
                  if (6'h1f == _T_288) begin
                    mem_31 <= _GEN_27;
                  end else begin
                    if (6'h1f == _T_283) begin
                      mem_31 <= _GEN_26;
                    end else begin
                      if (6'h1f == _T_278) begin
                        mem_31 <= _GEN_25;
                      end else begin
                        if (6'h1f == _T_273) begin
                          mem_31 <= _GEN_24;
                        end else begin
                          if (6'h1f == _T_268) begin
                            mem_31 <= _GEN_23;
                          end else begin
                            if (6'h1f == _T_263) begin
                              mem_31 <= _GEN_22;
                            end else begin
                              if (6'h1f == _T_258) begin
                                mem_31 <= _GEN_21;
                              end else begin
                                if (6'h1f == _T_253) begin
                                  mem_31 <= _GEN_20;
                                end else begin
                                  if (6'h1f == _T_248) begin
                                    mem_31 <= _GEN_19;
                                  end else begin
                                    if (6'h1f == _T_243) begin
                                      mem_31 <= _GEN_18;
                                    end else begin
                                      if (6'h1f == _T_238) begin
                                        mem_31 <= _GEN_17;
                                      end else begin
                                        if (6'h1f == _T_233) begin
                                          mem_31 <= _GEN_16;
                                        end else begin
                                          if (6'h1f == _T_228) begin
                                            mem_31 <= _GEN_15;
                                          end else begin
                                            if (6'h1f == _T_223) begin
                                              mem_31 <= _GEN_14;
                                            end else begin
                                              if (6'h1f == _T_218) begin
                                                mem_31 <= _GEN_13;
                                              end else begin
                                                if (6'h1f == _T_213) begin
                                                  mem_31 <= _GEN_12;
                                                end else begin
                                                  if (6'h1f == _T_208) begin
                                                    mem_31 <= _GEN_11;
                                                  end else begin
                                                    if (6'h1f == _T_203) begin
                                                      mem_31 <= _GEN_10;
                                                    end else begin
                                                      if (6'h1f == _T_198) begin
                                                        mem_31 <= _GEN_9;
                                                      end else begin
                                                        if (6'h1f == _T_193) begin
                                                          mem_31 <= _GEN_8;
                                                        end else begin
                                                          if (6'h1f == _T_188) begin
                                                            mem_31 <= _GEN_7;
                                                          end else begin
                                                            if (6'h1f == _T_183) begin
                                                              mem_31 <= _GEN_6;
                                                            end else begin
                                                              if (6'h1f == _T_178) begin
                                                                mem_31 <= _GEN_5;
                                                              end else begin
                                                                if (6'h1f == _T_173) begin
                                                                  mem_31 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h1f == _T_168) begin
                                                                    mem_31 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h1f == _T_163) begin
                                                                      mem_31 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h1f == _T_158) begin
                                                                        mem_31 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h1f == _T_153) begin
                                                                          mem_31 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h1f == _T_308) begin
          mem_31 <= _GEN_31;
        end else begin
          if (6'h1f == _T_303) begin
            mem_31 <= _GEN_30;
          end else begin
            if (6'h1f == _T_298) begin
              mem_31 <= _GEN_29;
            end else begin
              if (6'h1f == _T_293) begin
                mem_31 <= _GEN_28;
              end else begin
                if (6'h1f == _T_288) begin
                  mem_31 <= _GEN_27;
                end else begin
                  if (6'h1f == _T_283) begin
                    mem_31 <= _GEN_26;
                  end else begin
                    if (6'h1f == _T_278) begin
                      mem_31 <= _GEN_25;
                    end else begin
                      if (6'h1f == _T_273) begin
                        mem_31 <= _GEN_24;
                      end else begin
                        if (6'h1f == _T_268) begin
                          mem_31 <= _GEN_23;
                        end else begin
                          if (6'h1f == _T_263) begin
                            mem_31 <= _GEN_22;
                          end else begin
                            if (6'h1f == _T_258) begin
                              mem_31 <= _GEN_21;
                            end else begin
                              if (6'h1f == _T_253) begin
                                mem_31 <= _GEN_20;
                              end else begin
                                if (6'h1f == _T_248) begin
                                  mem_31 <= _GEN_19;
                                end else begin
                                  if (6'h1f == _T_243) begin
                                    mem_31 <= _GEN_18;
                                  end else begin
                                    if (6'h1f == _T_238) begin
                                      mem_31 <= _GEN_17;
                                    end else begin
                                      if (6'h1f == _T_233) begin
                                        mem_31 <= _GEN_16;
                                      end else begin
                                        if (6'h1f == _T_228) begin
                                          mem_31 <= _GEN_15;
                                        end else begin
                                          if (6'h1f == _T_223) begin
                                            mem_31 <= _GEN_14;
                                          end else begin
                                            if (6'h1f == _T_218) begin
                                              mem_31 <= _GEN_13;
                                            end else begin
                                              if (6'h1f == _T_213) begin
                                                mem_31 <= _GEN_12;
                                              end else begin
                                                if (6'h1f == _T_208) begin
                                                  mem_31 <= _GEN_11;
                                                end else begin
                                                  if (6'h1f == _T_203) begin
                                                    mem_31 <= _GEN_10;
                                                  end else begin
                                                    if (6'h1f == _T_198) begin
                                                      mem_31 <= _GEN_9;
                                                    end else begin
                                                      if (6'h1f == _T_193) begin
                                                        mem_31 <= _GEN_8;
                                                      end else begin
                                                        if (6'h1f == _T_188) begin
                                                          mem_31 <= _GEN_7;
                                                        end else begin
                                                          if (6'h1f == _T_183) begin
                                                            mem_31 <= _GEN_6;
                                                          end else begin
                                                            if (6'h1f == _T_178) begin
                                                              mem_31 <= _GEN_5;
                                                            end else begin
                                                              if (6'h1f == _T_173) begin
                                                                mem_31 <= _GEN_4;
                                                              end else begin
                                                                if (6'h1f == _T_168) begin
                                                                  mem_31 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h1f == _T_163) begin
                                                                    mem_31 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h1f == _T_158) begin
                                                                      mem_31 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h1f == _T_153) begin
                                                                        mem_31 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h20 == wPos) begin
            mem_32 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h20 == _T_308) begin
                mem_32 <= _GEN_31;
              end else begin
                if (6'h20 == _T_303) begin
                  mem_32 <= _GEN_30;
                end else begin
                  if (6'h20 == _T_298) begin
                    mem_32 <= _GEN_29;
                  end else begin
                    if (6'h20 == _T_293) begin
                      mem_32 <= _GEN_28;
                    end else begin
                      if (6'h20 == _T_288) begin
                        mem_32 <= _GEN_27;
                      end else begin
                        if (6'h20 == _T_283) begin
                          mem_32 <= _GEN_26;
                        end else begin
                          if (6'h20 == _T_278) begin
                            mem_32 <= _GEN_25;
                          end else begin
                            if (6'h20 == _T_273) begin
                              mem_32 <= _GEN_24;
                            end else begin
                              if (6'h20 == _T_268) begin
                                mem_32 <= _GEN_23;
                              end else begin
                                if (6'h20 == _T_263) begin
                                  mem_32 <= _GEN_22;
                                end else begin
                                  if (6'h20 == _T_258) begin
                                    mem_32 <= _GEN_21;
                                  end else begin
                                    if (6'h20 == _T_253) begin
                                      mem_32 <= _GEN_20;
                                    end else begin
                                      if (6'h20 == _T_248) begin
                                        mem_32 <= _GEN_19;
                                      end else begin
                                        if (6'h20 == _T_243) begin
                                          mem_32 <= _GEN_18;
                                        end else begin
                                          if (6'h20 == _T_238) begin
                                            mem_32 <= _GEN_17;
                                          end else begin
                                            if (6'h20 == _T_233) begin
                                              mem_32 <= _GEN_16;
                                            end else begin
                                              if (6'h20 == _T_228) begin
                                                mem_32 <= _GEN_15;
                                              end else begin
                                                if (6'h20 == _T_223) begin
                                                  mem_32 <= _GEN_14;
                                                end else begin
                                                  if (6'h20 == _T_218) begin
                                                    mem_32 <= _GEN_13;
                                                  end else begin
                                                    if (6'h20 == _T_213) begin
                                                      mem_32 <= _GEN_12;
                                                    end else begin
                                                      if (6'h20 == _T_208) begin
                                                        mem_32 <= _GEN_11;
                                                      end else begin
                                                        if (6'h20 == _T_203) begin
                                                          mem_32 <= _GEN_10;
                                                        end else begin
                                                          if (6'h20 == _T_198) begin
                                                            mem_32 <= _GEN_9;
                                                          end else begin
                                                            if (6'h20 == _T_193) begin
                                                              mem_32 <= _GEN_8;
                                                            end else begin
                                                              if (6'h20 == _T_188) begin
                                                                mem_32 <= _GEN_7;
                                                              end else begin
                                                                if (6'h20 == _T_183) begin
                                                                  mem_32 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h20 == _T_178) begin
                                                                    mem_32 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h20 == _T_173) begin
                                                                      mem_32 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h20 == _T_168) begin
                                                                        mem_32 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h20 == _T_163) begin
                                                                          mem_32 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h20 == _T_158) begin
                                                                            mem_32 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h20 == _T_153) begin
                                                                              mem_32 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h20 == _T_308) begin
              mem_32 <= _GEN_31;
            end else begin
              if (6'h20 == _T_303) begin
                mem_32 <= _GEN_30;
              end else begin
                if (6'h20 == _T_298) begin
                  mem_32 <= _GEN_29;
                end else begin
                  if (6'h20 == _T_293) begin
                    mem_32 <= _GEN_28;
                  end else begin
                    if (6'h20 == _T_288) begin
                      mem_32 <= _GEN_27;
                    end else begin
                      if (6'h20 == _T_283) begin
                        mem_32 <= _GEN_26;
                      end else begin
                        if (6'h20 == _T_278) begin
                          mem_32 <= _GEN_25;
                        end else begin
                          if (6'h20 == _T_273) begin
                            mem_32 <= _GEN_24;
                          end else begin
                            if (6'h20 == _T_268) begin
                              mem_32 <= _GEN_23;
                            end else begin
                              if (6'h20 == _T_263) begin
                                mem_32 <= _GEN_22;
                              end else begin
                                if (6'h20 == _T_258) begin
                                  mem_32 <= _GEN_21;
                                end else begin
                                  if (6'h20 == _T_253) begin
                                    mem_32 <= _GEN_20;
                                  end else begin
                                    if (6'h20 == _T_248) begin
                                      mem_32 <= _GEN_19;
                                    end else begin
                                      if (6'h20 == _T_243) begin
                                        mem_32 <= _GEN_18;
                                      end else begin
                                        if (6'h20 == _T_238) begin
                                          mem_32 <= _GEN_17;
                                        end else begin
                                          if (6'h20 == _T_233) begin
                                            mem_32 <= _GEN_16;
                                          end else begin
                                            if (6'h20 == _T_228) begin
                                              mem_32 <= _GEN_15;
                                            end else begin
                                              if (6'h20 == _T_223) begin
                                                mem_32 <= _GEN_14;
                                              end else begin
                                                if (6'h20 == _T_218) begin
                                                  mem_32 <= _GEN_13;
                                                end else begin
                                                  if (6'h20 == _T_213) begin
                                                    mem_32 <= _GEN_12;
                                                  end else begin
                                                    if (6'h20 == _T_208) begin
                                                      mem_32 <= _GEN_11;
                                                    end else begin
                                                      if (6'h20 == _T_203) begin
                                                        mem_32 <= _GEN_10;
                                                      end else begin
                                                        if (6'h20 == _T_198) begin
                                                          mem_32 <= _GEN_9;
                                                        end else begin
                                                          if (6'h20 == _T_193) begin
                                                            mem_32 <= _GEN_8;
                                                          end else begin
                                                            if (6'h20 == _T_188) begin
                                                              mem_32 <= _GEN_7;
                                                            end else begin
                                                              if (6'h20 == _T_183) begin
                                                                mem_32 <= _GEN_6;
                                                              end else begin
                                                                if (6'h20 == _T_178) begin
                                                                  mem_32 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h20 == _T_173) begin
                                                                    mem_32 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h20 == _T_168) begin
                                                                      mem_32 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h20 == _T_163) begin
                                                                        mem_32 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h20 == _T_158) begin
                                                                          mem_32 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h20 == _T_153) begin
                                                                            mem_32 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h20 == _T_308) begin
            mem_32 <= _GEN_31;
          end else begin
            if (6'h20 == _T_303) begin
              mem_32 <= _GEN_30;
            end else begin
              if (6'h20 == _T_298) begin
                mem_32 <= _GEN_29;
              end else begin
                if (6'h20 == _T_293) begin
                  mem_32 <= _GEN_28;
                end else begin
                  if (6'h20 == _T_288) begin
                    mem_32 <= _GEN_27;
                  end else begin
                    if (6'h20 == _T_283) begin
                      mem_32 <= _GEN_26;
                    end else begin
                      if (6'h20 == _T_278) begin
                        mem_32 <= _GEN_25;
                      end else begin
                        if (6'h20 == _T_273) begin
                          mem_32 <= _GEN_24;
                        end else begin
                          if (6'h20 == _T_268) begin
                            mem_32 <= _GEN_23;
                          end else begin
                            if (6'h20 == _T_263) begin
                              mem_32 <= _GEN_22;
                            end else begin
                              if (6'h20 == _T_258) begin
                                mem_32 <= _GEN_21;
                              end else begin
                                if (6'h20 == _T_253) begin
                                  mem_32 <= _GEN_20;
                                end else begin
                                  if (6'h20 == _T_248) begin
                                    mem_32 <= _GEN_19;
                                  end else begin
                                    if (6'h20 == _T_243) begin
                                      mem_32 <= _GEN_18;
                                    end else begin
                                      if (6'h20 == _T_238) begin
                                        mem_32 <= _GEN_17;
                                      end else begin
                                        if (6'h20 == _T_233) begin
                                          mem_32 <= _GEN_16;
                                        end else begin
                                          if (6'h20 == _T_228) begin
                                            mem_32 <= _GEN_15;
                                          end else begin
                                            if (6'h20 == _T_223) begin
                                              mem_32 <= _GEN_14;
                                            end else begin
                                              if (6'h20 == _T_218) begin
                                                mem_32 <= _GEN_13;
                                              end else begin
                                                if (6'h20 == _T_213) begin
                                                  mem_32 <= _GEN_12;
                                                end else begin
                                                  if (6'h20 == _T_208) begin
                                                    mem_32 <= _GEN_11;
                                                  end else begin
                                                    if (6'h20 == _T_203) begin
                                                      mem_32 <= _GEN_10;
                                                    end else begin
                                                      if (6'h20 == _T_198) begin
                                                        mem_32 <= _GEN_9;
                                                      end else begin
                                                        if (6'h20 == _T_193) begin
                                                          mem_32 <= _GEN_8;
                                                        end else begin
                                                          if (6'h20 == _T_188) begin
                                                            mem_32 <= _GEN_7;
                                                          end else begin
                                                            if (6'h20 == _T_183) begin
                                                              mem_32 <= _GEN_6;
                                                            end else begin
                                                              if (6'h20 == _T_178) begin
                                                                mem_32 <= _GEN_5;
                                                              end else begin
                                                                if (6'h20 == _T_173) begin
                                                                  mem_32 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h20 == _T_168) begin
                                                                    mem_32 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h20 == _T_163) begin
                                                                      mem_32 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h20 == _T_158) begin
                                                                        mem_32 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h20 == _T_153) begin
                                                                          mem_32 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h20 == _T_308) begin
          mem_32 <= _GEN_31;
        end else begin
          if (6'h20 == _T_303) begin
            mem_32 <= _GEN_30;
          end else begin
            if (6'h20 == _T_298) begin
              mem_32 <= _GEN_29;
            end else begin
              if (6'h20 == _T_293) begin
                mem_32 <= _GEN_28;
              end else begin
                if (6'h20 == _T_288) begin
                  mem_32 <= _GEN_27;
                end else begin
                  if (6'h20 == _T_283) begin
                    mem_32 <= _GEN_26;
                  end else begin
                    if (6'h20 == _T_278) begin
                      mem_32 <= _GEN_25;
                    end else begin
                      if (6'h20 == _T_273) begin
                        mem_32 <= _GEN_24;
                      end else begin
                        if (6'h20 == _T_268) begin
                          mem_32 <= _GEN_23;
                        end else begin
                          if (6'h20 == _T_263) begin
                            mem_32 <= _GEN_22;
                          end else begin
                            if (6'h20 == _T_258) begin
                              mem_32 <= _GEN_21;
                            end else begin
                              if (6'h20 == _T_253) begin
                                mem_32 <= _GEN_20;
                              end else begin
                                if (6'h20 == _T_248) begin
                                  mem_32 <= _GEN_19;
                                end else begin
                                  if (6'h20 == _T_243) begin
                                    mem_32 <= _GEN_18;
                                  end else begin
                                    if (6'h20 == _T_238) begin
                                      mem_32 <= _GEN_17;
                                    end else begin
                                      if (6'h20 == _T_233) begin
                                        mem_32 <= _GEN_16;
                                      end else begin
                                        if (6'h20 == _T_228) begin
                                          mem_32 <= _GEN_15;
                                        end else begin
                                          if (6'h20 == _T_223) begin
                                            mem_32 <= _GEN_14;
                                          end else begin
                                            if (6'h20 == _T_218) begin
                                              mem_32 <= _GEN_13;
                                            end else begin
                                              if (6'h20 == _T_213) begin
                                                mem_32 <= _GEN_12;
                                              end else begin
                                                if (6'h20 == _T_208) begin
                                                  mem_32 <= _GEN_11;
                                                end else begin
                                                  if (6'h20 == _T_203) begin
                                                    mem_32 <= _GEN_10;
                                                  end else begin
                                                    if (6'h20 == _T_198) begin
                                                      mem_32 <= _GEN_9;
                                                    end else begin
                                                      if (6'h20 == _T_193) begin
                                                        mem_32 <= _GEN_8;
                                                      end else begin
                                                        if (6'h20 == _T_188) begin
                                                          mem_32 <= _GEN_7;
                                                        end else begin
                                                          if (6'h20 == _T_183) begin
                                                            mem_32 <= _GEN_6;
                                                          end else begin
                                                            if (6'h20 == _T_178) begin
                                                              mem_32 <= _GEN_5;
                                                            end else begin
                                                              if (6'h20 == _T_173) begin
                                                                mem_32 <= _GEN_4;
                                                              end else begin
                                                                if (6'h20 == _T_168) begin
                                                                  mem_32 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h20 == _T_163) begin
                                                                    mem_32 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h20 == _T_158) begin
                                                                      mem_32 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h20 == _T_153) begin
                                                                        mem_32 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h21 == wPos) begin
            mem_33 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h21 == _T_308) begin
                mem_33 <= _GEN_31;
              end else begin
                if (6'h21 == _T_303) begin
                  mem_33 <= _GEN_30;
                end else begin
                  if (6'h21 == _T_298) begin
                    mem_33 <= _GEN_29;
                  end else begin
                    if (6'h21 == _T_293) begin
                      mem_33 <= _GEN_28;
                    end else begin
                      if (6'h21 == _T_288) begin
                        mem_33 <= _GEN_27;
                      end else begin
                        if (6'h21 == _T_283) begin
                          mem_33 <= _GEN_26;
                        end else begin
                          if (6'h21 == _T_278) begin
                            mem_33 <= _GEN_25;
                          end else begin
                            if (6'h21 == _T_273) begin
                              mem_33 <= _GEN_24;
                            end else begin
                              if (6'h21 == _T_268) begin
                                mem_33 <= _GEN_23;
                              end else begin
                                if (6'h21 == _T_263) begin
                                  mem_33 <= _GEN_22;
                                end else begin
                                  if (6'h21 == _T_258) begin
                                    mem_33 <= _GEN_21;
                                  end else begin
                                    if (6'h21 == _T_253) begin
                                      mem_33 <= _GEN_20;
                                    end else begin
                                      if (6'h21 == _T_248) begin
                                        mem_33 <= _GEN_19;
                                      end else begin
                                        if (6'h21 == _T_243) begin
                                          mem_33 <= _GEN_18;
                                        end else begin
                                          if (6'h21 == _T_238) begin
                                            mem_33 <= _GEN_17;
                                          end else begin
                                            if (6'h21 == _T_233) begin
                                              mem_33 <= _GEN_16;
                                            end else begin
                                              if (6'h21 == _T_228) begin
                                                mem_33 <= _GEN_15;
                                              end else begin
                                                if (6'h21 == _T_223) begin
                                                  mem_33 <= _GEN_14;
                                                end else begin
                                                  if (6'h21 == _T_218) begin
                                                    mem_33 <= _GEN_13;
                                                  end else begin
                                                    if (6'h21 == _T_213) begin
                                                      mem_33 <= _GEN_12;
                                                    end else begin
                                                      if (6'h21 == _T_208) begin
                                                        mem_33 <= _GEN_11;
                                                      end else begin
                                                        if (6'h21 == _T_203) begin
                                                          mem_33 <= _GEN_10;
                                                        end else begin
                                                          if (6'h21 == _T_198) begin
                                                            mem_33 <= _GEN_9;
                                                          end else begin
                                                            if (6'h21 == _T_193) begin
                                                              mem_33 <= _GEN_8;
                                                            end else begin
                                                              if (6'h21 == _T_188) begin
                                                                mem_33 <= _GEN_7;
                                                              end else begin
                                                                if (6'h21 == _T_183) begin
                                                                  mem_33 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h21 == _T_178) begin
                                                                    mem_33 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h21 == _T_173) begin
                                                                      mem_33 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h21 == _T_168) begin
                                                                        mem_33 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h21 == _T_163) begin
                                                                          mem_33 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h21 == _T_158) begin
                                                                            mem_33 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h21 == _T_153) begin
                                                                              mem_33 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h21 == _T_308) begin
              mem_33 <= _GEN_31;
            end else begin
              if (6'h21 == _T_303) begin
                mem_33 <= _GEN_30;
              end else begin
                if (6'h21 == _T_298) begin
                  mem_33 <= _GEN_29;
                end else begin
                  if (6'h21 == _T_293) begin
                    mem_33 <= _GEN_28;
                  end else begin
                    if (6'h21 == _T_288) begin
                      mem_33 <= _GEN_27;
                    end else begin
                      if (6'h21 == _T_283) begin
                        mem_33 <= _GEN_26;
                      end else begin
                        if (6'h21 == _T_278) begin
                          mem_33 <= _GEN_25;
                        end else begin
                          if (6'h21 == _T_273) begin
                            mem_33 <= _GEN_24;
                          end else begin
                            if (6'h21 == _T_268) begin
                              mem_33 <= _GEN_23;
                            end else begin
                              if (6'h21 == _T_263) begin
                                mem_33 <= _GEN_22;
                              end else begin
                                if (6'h21 == _T_258) begin
                                  mem_33 <= _GEN_21;
                                end else begin
                                  if (6'h21 == _T_253) begin
                                    mem_33 <= _GEN_20;
                                  end else begin
                                    if (6'h21 == _T_248) begin
                                      mem_33 <= _GEN_19;
                                    end else begin
                                      if (6'h21 == _T_243) begin
                                        mem_33 <= _GEN_18;
                                      end else begin
                                        if (6'h21 == _T_238) begin
                                          mem_33 <= _GEN_17;
                                        end else begin
                                          if (6'h21 == _T_233) begin
                                            mem_33 <= _GEN_16;
                                          end else begin
                                            if (6'h21 == _T_228) begin
                                              mem_33 <= _GEN_15;
                                            end else begin
                                              if (6'h21 == _T_223) begin
                                                mem_33 <= _GEN_14;
                                              end else begin
                                                if (6'h21 == _T_218) begin
                                                  mem_33 <= _GEN_13;
                                                end else begin
                                                  if (6'h21 == _T_213) begin
                                                    mem_33 <= _GEN_12;
                                                  end else begin
                                                    if (6'h21 == _T_208) begin
                                                      mem_33 <= _GEN_11;
                                                    end else begin
                                                      if (6'h21 == _T_203) begin
                                                        mem_33 <= _GEN_10;
                                                      end else begin
                                                        if (6'h21 == _T_198) begin
                                                          mem_33 <= _GEN_9;
                                                        end else begin
                                                          if (6'h21 == _T_193) begin
                                                            mem_33 <= _GEN_8;
                                                          end else begin
                                                            if (6'h21 == _T_188) begin
                                                              mem_33 <= _GEN_7;
                                                            end else begin
                                                              if (6'h21 == _T_183) begin
                                                                mem_33 <= _GEN_6;
                                                              end else begin
                                                                if (6'h21 == _T_178) begin
                                                                  mem_33 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h21 == _T_173) begin
                                                                    mem_33 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h21 == _T_168) begin
                                                                      mem_33 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h21 == _T_163) begin
                                                                        mem_33 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h21 == _T_158) begin
                                                                          mem_33 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h21 == _T_153) begin
                                                                            mem_33 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h21 == _T_308) begin
            mem_33 <= _GEN_31;
          end else begin
            if (6'h21 == _T_303) begin
              mem_33 <= _GEN_30;
            end else begin
              if (6'h21 == _T_298) begin
                mem_33 <= _GEN_29;
              end else begin
                if (6'h21 == _T_293) begin
                  mem_33 <= _GEN_28;
                end else begin
                  if (6'h21 == _T_288) begin
                    mem_33 <= _GEN_27;
                  end else begin
                    if (6'h21 == _T_283) begin
                      mem_33 <= _GEN_26;
                    end else begin
                      if (6'h21 == _T_278) begin
                        mem_33 <= _GEN_25;
                      end else begin
                        if (6'h21 == _T_273) begin
                          mem_33 <= _GEN_24;
                        end else begin
                          if (6'h21 == _T_268) begin
                            mem_33 <= _GEN_23;
                          end else begin
                            if (6'h21 == _T_263) begin
                              mem_33 <= _GEN_22;
                            end else begin
                              if (6'h21 == _T_258) begin
                                mem_33 <= _GEN_21;
                              end else begin
                                if (6'h21 == _T_253) begin
                                  mem_33 <= _GEN_20;
                                end else begin
                                  if (6'h21 == _T_248) begin
                                    mem_33 <= _GEN_19;
                                  end else begin
                                    if (6'h21 == _T_243) begin
                                      mem_33 <= _GEN_18;
                                    end else begin
                                      if (6'h21 == _T_238) begin
                                        mem_33 <= _GEN_17;
                                      end else begin
                                        if (6'h21 == _T_233) begin
                                          mem_33 <= _GEN_16;
                                        end else begin
                                          if (6'h21 == _T_228) begin
                                            mem_33 <= _GEN_15;
                                          end else begin
                                            if (6'h21 == _T_223) begin
                                              mem_33 <= _GEN_14;
                                            end else begin
                                              if (6'h21 == _T_218) begin
                                                mem_33 <= _GEN_13;
                                              end else begin
                                                if (6'h21 == _T_213) begin
                                                  mem_33 <= _GEN_12;
                                                end else begin
                                                  if (6'h21 == _T_208) begin
                                                    mem_33 <= _GEN_11;
                                                  end else begin
                                                    if (6'h21 == _T_203) begin
                                                      mem_33 <= _GEN_10;
                                                    end else begin
                                                      if (6'h21 == _T_198) begin
                                                        mem_33 <= _GEN_9;
                                                      end else begin
                                                        if (6'h21 == _T_193) begin
                                                          mem_33 <= _GEN_8;
                                                        end else begin
                                                          if (6'h21 == _T_188) begin
                                                            mem_33 <= _GEN_7;
                                                          end else begin
                                                            if (6'h21 == _T_183) begin
                                                              mem_33 <= _GEN_6;
                                                            end else begin
                                                              if (6'h21 == _T_178) begin
                                                                mem_33 <= _GEN_5;
                                                              end else begin
                                                                if (6'h21 == _T_173) begin
                                                                  mem_33 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h21 == _T_168) begin
                                                                    mem_33 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h21 == _T_163) begin
                                                                      mem_33 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h21 == _T_158) begin
                                                                        mem_33 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h21 == _T_153) begin
                                                                          mem_33 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h21 == _T_308) begin
          mem_33 <= _GEN_31;
        end else begin
          if (6'h21 == _T_303) begin
            mem_33 <= _GEN_30;
          end else begin
            if (6'h21 == _T_298) begin
              mem_33 <= _GEN_29;
            end else begin
              if (6'h21 == _T_293) begin
                mem_33 <= _GEN_28;
              end else begin
                if (6'h21 == _T_288) begin
                  mem_33 <= _GEN_27;
                end else begin
                  if (6'h21 == _T_283) begin
                    mem_33 <= _GEN_26;
                  end else begin
                    if (6'h21 == _T_278) begin
                      mem_33 <= _GEN_25;
                    end else begin
                      if (6'h21 == _T_273) begin
                        mem_33 <= _GEN_24;
                      end else begin
                        if (6'h21 == _T_268) begin
                          mem_33 <= _GEN_23;
                        end else begin
                          if (6'h21 == _T_263) begin
                            mem_33 <= _GEN_22;
                          end else begin
                            if (6'h21 == _T_258) begin
                              mem_33 <= _GEN_21;
                            end else begin
                              if (6'h21 == _T_253) begin
                                mem_33 <= _GEN_20;
                              end else begin
                                if (6'h21 == _T_248) begin
                                  mem_33 <= _GEN_19;
                                end else begin
                                  if (6'h21 == _T_243) begin
                                    mem_33 <= _GEN_18;
                                  end else begin
                                    if (6'h21 == _T_238) begin
                                      mem_33 <= _GEN_17;
                                    end else begin
                                      if (6'h21 == _T_233) begin
                                        mem_33 <= _GEN_16;
                                      end else begin
                                        if (6'h21 == _T_228) begin
                                          mem_33 <= _GEN_15;
                                        end else begin
                                          if (6'h21 == _T_223) begin
                                            mem_33 <= _GEN_14;
                                          end else begin
                                            if (6'h21 == _T_218) begin
                                              mem_33 <= _GEN_13;
                                            end else begin
                                              if (6'h21 == _T_213) begin
                                                mem_33 <= _GEN_12;
                                              end else begin
                                                if (6'h21 == _T_208) begin
                                                  mem_33 <= _GEN_11;
                                                end else begin
                                                  if (6'h21 == _T_203) begin
                                                    mem_33 <= _GEN_10;
                                                  end else begin
                                                    if (6'h21 == _T_198) begin
                                                      mem_33 <= _GEN_9;
                                                    end else begin
                                                      if (6'h21 == _T_193) begin
                                                        mem_33 <= _GEN_8;
                                                      end else begin
                                                        if (6'h21 == _T_188) begin
                                                          mem_33 <= _GEN_7;
                                                        end else begin
                                                          if (6'h21 == _T_183) begin
                                                            mem_33 <= _GEN_6;
                                                          end else begin
                                                            if (6'h21 == _T_178) begin
                                                              mem_33 <= _GEN_5;
                                                            end else begin
                                                              if (6'h21 == _T_173) begin
                                                                mem_33 <= _GEN_4;
                                                              end else begin
                                                                if (6'h21 == _T_168) begin
                                                                  mem_33 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h21 == _T_163) begin
                                                                    mem_33 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h21 == _T_158) begin
                                                                      mem_33 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h21 == _T_153) begin
                                                                        mem_33 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h22 == wPos) begin
            mem_34 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h22 == _T_308) begin
                mem_34 <= _GEN_31;
              end else begin
                if (6'h22 == _T_303) begin
                  mem_34 <= _GEN_30;
                end else begin
                  if (6'h22 == _T_298) begin
                    mem_34 <= _GEN_29;
                  end else begin
                    if (6'h22 == _T_293) begin
                      mem_34 <= _GEN_28;
                    end else begin
                      if (6'h22 == _T_288) begin
                        mem_34 <= _GEN_27;
                      end else begin
                        if (6'h22 == _T_283) begin
                          mem_34 <= _GEN_26;
                        end else begin
                          if (6'h22 == _T_278) begin
                            mem_34 <= _GEN_25;
                          end else begin
                            if (6'h22 == _T_273) begin
                              mem_34 <= _GEN_24;
                            end else begin
                              if (6'h22 == _T_268) begin
                                mem_34 <= _GEN_23;
                              end else begin
                                if (6'h22 == _T_263) begin
                                  mem_34 <= _GEN_22;
                                end else begin
                                  if (6'h22 == _T_258) begin
                                    mem_34 <= _GEN_21;
                                  end else begin
                                    if (6'h22 == _T_253) begin
                                      mem_34 <= _GEN_20;
                                    end else begin
                                      if (6'h22 == _T_248) begin
                                        mem_34 <= _GEN_19;
                                      end else begin
                                        if (6'h22 == _T_243) begin
                                          mem_34 <= _GEN_18;
                                        end else begin
                                          if (6'h22 == _T_238) begin
                                            mem_34 <= _GEN_17;
                                          end else begin
                                            if (6'h22 == _T_233) begin
                                              mem_34 <= _GEN_16;
                                            end else begin
                                              if (6'h22 == _T_228) begin
                                                mem_34 <= _GEN_15;
                                              end else begin
                                                if (6'h22 == _T_223) begin
                                                  mem_34 <= _GEN_14;
                                                end else begin
                                                  if (6'h22 == _T_218) begin
                                                    mem_34 <= _GEN_13;
                                                  end else begin
                                                    if (6'h22 == _T_213) begin
                                                      mem_34 <= _GEN_12;
                                                    end else begin
                                                      if (6'h22 == _T_208) begin
                                                        mem_34 <= _GEN_11;
                                                      end else begin
                                                        if (6'h22 == _T_203) begin
                                                          mem_34 <= _GEN_10;
                                                        end else begin
                                                          if (6'h22 == _T_198) begin
                                                            mem_34 <= _GEN_9;
                                                          end else begin
                                                            if (6'h22 == _T_193) begin
                                                              mem_34 <= _GEN_8;
                                                            end else begin
                                                              if (6'h22 == _T_188) begin
                                                                mem_34 <= _GEN_7;
                                                              end else begin
                                                                if (6'h22 == _T_183) begin
                                                                  mem_34 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h22 == _T_178) begin
                                                                    mem_34 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h22 == _T_173) begin
                                                                      mem_34 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h22 == _T_168) begin
                                                                        mem_34 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h22 == _T_163) begin
                                                                          mem_34 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h22 == _T_158) begin
                                                                            mem_34 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h22 == _T_153) begin
                                                                              mem_34 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h22 == _T_308) begin
              mem_34 <= _GEN_31;
            end else begin
              if (6'h22 == _T_303) begin
                mem_34 <= _GEN_30;
              end else begin
                if (6'h22 == _T_298) begin
                  mem_34 <= _GEN_29;
                end else begin
                  if (6'h22 == _T_293) begin
                    mem_34 <= _GEN_28;
                  end else begin
                    if (6'h22 == _T_288) begin
                      mem_34 <= _GEN_27;
                    end else begin
                      if (6'h22 == _T_283) begin
                        mem_34 <= _GEN_26;
                      end else begin
                        if (6'h22 == _T_278) begin
                          mem_34 <= _GEN_25;
                        end else begin
                          if (6'h22 == _T_273) begin
                            mem_34 <= _GEN_24;
                          end else begin
                            if (6'h22 == _T_268) begin
                              mem_34 <= _GEN_23;
                            end else begin
                              if (6'h22 == _T_263) begin
                                mem_34 <= _GEN_22;
                              end else begin
                                if (6'h22 == _T_258) begin
                                  mem_34 <= _GEN_21;
                                end else begin
                                  if (6'h22 == _T_253) begin
                                    mem_34 <= _GEN_20;
                                  end else begin
                                    if (6'h22 == _T_248) begin
                                      mem_34 <= _GEN_19;
                                    end else begin
                                      if (6'h22 == _T_243) begin
                                        mem_34 <= _GEN_18;
                                      end else begin
                                        if (6'h22 == _T_238) begin
                                          mem_34 <= _GEN_17;
                                        end else begin
                                          if (6'h22 == _T_233) begin
                                            mem_34 <= _GEN_16;
                                          end else begin
                                            if (6'h22 == _T_228) begin
                                              mem_34 <= _GEN_15;
                                            end else begin
                                              if (6'h22 == _T_223) begin
                                                mem_34 <= _GEN_14;
                                              end else begin
                                                if (6'h22 == _T_218) begin
                                                  mem_34 <= _GEN_13;
                                                end else begin
                                                  if (6'h22 == _T_213) begin
                                                    mem_34 <= _GEN_12;
                                                  end else begin
                                                    if (6'h22 == _T_208) begin
                                                      mem_34 <= _GEN_11;
                                                    end else begin
                                                      if (6'h22 == _T_203) begin
                                                        mem_34 <= _GEN_10;
                                                      end else begin
                                                        if (6'h22 == _T_198) begin
                                                          mem_34 <= _GEN_9;
                                                        end else begin
                                                          if (6'h22 == _T_193) begin
                                                            mem_34 <= _GEN_8;
                                                          end else begin
                                                            if (6'h22 == _T_188) begin
                                                              mem_34 <= _GEN_7;
                                                            end else begin
                                                              if (6'h22 == _T_183) begin
                                                                mem_34 <= _GEN_6;
                                                              end else begin
                                                                if (6'h22 == _T_178) begin
                                                                  mem_34 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h22 == _T_173) begin
                                                                    mem_34 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h22 == _T_168) begin
                                                                      mem_34 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h22 == _T_163) begin
                                                                        mem_34 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h22 == _T_158) begin
                                                                          mem_34 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h22 == _T_153) begin
                                                                            mem_34 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h22 == _T_308) begin
            mem_34 <= _GEN_31;
          end else begin
            if (6'h22 == _T_303) begin
              mem_34 <= _GEN_30;
            end else begin
              if (6'h22 == _T_298) begin
                mem_34 <= _GEN_29;
              end else begin
                if (6'h22 == _T_293) begin
                  mem_34 <= _GEN_28;
                end else begin
                  if (6'h22 == _T_288) begin
                    mem_34 <= _GEN_27;
                  end else begin
                    if (6'h22 == _T_283) begin
                      mem_34 <= _GEN_26;
                    end else begin
                      if (6'h22 == _T_278) begin
                        mem_34 <= _GEN_25;
                      end else begin
                        if (6'h22 == _T_273) begin
                          mem_34 <= _GEN_24;
                        end else begin
                          if (6'h22 == _T_268) begin
                            mem_34 <= _GEN_23;
                          end else begin
                            if (6'h22 == _T_263) begin
                              mem_34 <= _GEN_22;
                            end else begin
                              if (6'h22 == _T_258) begin
                                mem_34 <= _GEN_21;
                              end else begin
                                if (6'h22 == _T_253) begin
                                  mem_34 <= _GEN_20;
                                end else begin
                                  if (6'h22 == _T_248) begin
                                    mem_34 <= _GEN_19;
                                  end else begin
                                    if (6'h22 == _T_243) begin
                                      mem_34 <= _GEN_18;
                                    end else begin
                                      if (6'h22 == _T_238) begin
                                        mem_34 <= _GEN_17;
                                      end else begin
                                        if (6'h22 == _T_233) begin
                                          mem_34 <= _GEN_16;
                                        end else begin
                                          if (6'h22 == _T_228) begin
                                            mem_34 <= _GEN_15;
                                          end else begin
                                            if (6'h22 == _T_223) begin
                                              mem_34 <= _GEN_14;
                                            end else begin
                                              if (6'h22 == _T_218) begin
                                                mem_34 <= _GEN_13;
                                              end else begin
                                                if (6'h22 == _T_213) begin
                                                  mem_34 <= _GEN_12;
                                                end else begin
                                                  if (6'h22 == _T_208) begin
                                                    mem_34 <= _GEN_11;
                                                  end else begin
                                                    if (6'h22 == _T_203) begin
                                                      mem_34 <= _GEN_10;
                                                    end else begin
                                                      if (6'h22 == _T_198) begin
                                                        mem_34 <= _GEN_9;
                                                      end else begin
                                                        if (6'h22 == _T_193) begin
                                                          mem_34 <= _GEN_8;
                                                        end else begin
                                                          if (6'h22 == _T_188) begin
                                                            mem_34 <= _GEN_7;
                                                          end else begin
                                                            if (6'h22 == _T_183) begin
                                                              mem_34 <= _GEN_6;
                                                            end else begin
                                                              if (6'h22 == _T_178) begin
                                                                mem_34 <= _GEN_5;
                                                              end else begin
                                                                if (6'h22 == _T_173) begin
                                                                  mem_34 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h22 == _T_168) begin
                                                                    mem_34 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h22 == _T_163) begin
                                                                      mem_34 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h22 == _T_158) begin
                                                                        mem_34 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h22 == _T_153) begin
                                                                          mem_34 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h22 == _T_308) begin
          mem_34 <= _GEN_31;
        end else begin
          if (6'h22 == _T_303) begin
            mem_34 <= _GEN_30;
          end else begin
            if (6'h22 == _T_298) begin
              mem_34 <= _GEN_29;
            end else begin
              if (6'h22 == _T_293) begin
                mem_34 <= _GEN_28;
              end else begin
                if (6'h22 == _T_288) begin
                  mem_34 <= _GEN_27;
                end else begin
                  if (6'h22 == _T_283) begin
                    mem_34 <= _GEN_26;
                  end else begin
                    if (6'h22 == _T_278) begin
                      mem_34 <= _GEN_25;
                    end else begin
                      if (6'h22 == _T_273) begin
                        mem_34 <= _GEN_24;
                      end else begin
                        if (6'h22 == _T_268) begin
                          mem_34 <= _GEN_23;
                        end else begin
                          if (6'h22 == _T_263) begin
                            mem_34 <= _GEN_22;
                          end else begin
                            if (6'h22 == _T_258) begin
                              mem_34 <= _GEN_21;
                            end else begin
                              if (6'h22 == _T_253) begin
                                mem_34 <= _GEN_20;
                              end else begin
                                if (6'h22 == _T_248) begin
                                  mem_34 <= _GEN_19;
                                end else begin
                                  if (6'h22 == _T_243) begin
                                    mem_34 <= _GEN_18;
                                  end else begin
                                    if (6'h22 == _T_238) begin
                                      mem_34 <= _GEN_17;
                                    end else begin
                                      if (6'h22 == _T_233) begin
                                        mem_34 <= _GEN_16;
                                      end else begin
                                        if (6'h22 == _T_228) begin
                                          mem_34 <= _GEN_15;
                                        end else begin
                                          if (6'h22 == _T_223) begin
                                            mem_34 <= _GEN_14;
                                          end else begin
                                            if (6'h22 == _T_218) begin
                                              mem_34 <= _GEN_13;
                                            end else begin
                                              if (6'h22 == _T_213) begin
                                                mem_34 <= _GEN_12;
                                              end else begin
                                                if (6'h22 == _T_208) begin
                                                  mem_34 <= _GEN_11;
                                                end else begin
                                                  if (6'h22 == _T_203) begin
                                                    mem_34 <= _GEN_10;
                                                  end else begin
                                                    if (6'h22 == _T_198) begin
                                                      mem_34 <= _GEN_9;
                                                    end else begin
                                                      if (6'h22 == _T_193) begin
                                                        mem_34 <= _GEN_8;
                                                      end else begin
                                                        if (6'h22 == _T_188) begin
                                                          mem_34 <= _GEN_7;
                                                        end else begin
                                                          if (6'h22 == _T_183) begin
                                                            mem_34 <= _GEN_6;
                                                          end else begin
                                                            if (6'h22 == _T_178) begin
                                                              mem_34 <= _GEN_5;
                                                            end else begin
                                                              if (6'h22 == _T_173) begin
                                                                mem_34 <= _GEN_4;
                                                              end else begin
                                                                if (6'h22 == _T_168) begin
                                                                  mem_34 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h22 == _T_163) begin
                                                                    mem_34 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h22 == _T_158) begin
                                                                      mem_34 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h22 == _T_153) begin
                                                                        mem_34 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h23 == wPos) begin
            mem_35 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h23 == _T_308) begin
                mem_35 <= _GEN_31;
              end else begin
                if (6'h23 == _T_303) begin
                  mem_35 <= _GEN_30;
                end else begin
                  if (6'h23 == _T_298) begin
                    mem_35 <= _GEN_29;
                  end else begin
                    if (6'h23 == _T_293) begin
                      mem_35 <= _GEN_28;
                    end else begin
                      if (6'h23 == _T_288) begin
                        mem_35 <= _GEN_27;
                      end else begin
                        if (6'h23 == _T_283) begin
                          mem_35 <= _GEN_26;
                        end else begin
                          if (6'h23 == _T_278) begin
                            mem_35 <= _GEN_25;
                          end else begin
                            if (6'h23 == _T_273) begin
                              mem_35 <= _GEN_24;
                            end else begin
                              if (6'h23 == _T_268) begin
                                mem_35 <= _GEN_23;
                              end else begin
                                if (6'h23 == _T_263) begin
                                  mem_35 <= _GEN_22;
                                end else begin
                                  if (6'h23 == _T_258) begin
                                    mem_35 <= _GEN_21;
                                  end else begin
                                    if (6'h23 == _T_253) begin
                                      mem_35 <= _GEN_20;
                                    end else begin
                                      if (6'h23 == _T_248) begin
                                        mem_35 <= _GEN_19;
                                      end else begin
                                        if (6'h23 == _T_243) begin
                                          mem_35 <= _GEN_18;
                                        end else begin
                                          if (6'h23 == _T_238) begin
                                            mem_35 <= _GEN_17;
                                          end else begin
                                            if (6'h23 == _T_233) begin
                                              mem_35 <= _GEN_16;
                                            end else begin
                                              if (6'h23 == _T_228) begin
                                                mem_35 <= _GEN_15;
                                              end else begin
                                                if (6'h23 == _T_223) begin
                                                  mem_35 <= _GEN_14;
                                                end else begin
                                                  if (6'h23 == _T_218) begin
                                                    mem_35 <= _GEN_13;
                                                  end else begin
                                                    if (6'h23 == _T_213) begin
                                                      mem_35 <= _GEN_12;
                                                    end else begin
                                                      if (6'h23 == _T_208) begin
                                                        mem_35 <= _GEN_11;
                                                      end else begin
                                                        if (6'h23 == _T_203) begin
                                                          mem_35 <= _GEN_10;
                                                        end else begin
                                                          if (6'h23 == _T_198) begin
                                                            mem_35 <= _GEN_9;
                                                          end else begin
                                                            if (6'h23 == _T_193) begin
                                                              mem_35 <= _GEN_8;
                                                            end else begin
                                                              if (6'h23 == _T_188) begin
                                                                mem_35 <= _GEN_7;
                                                              end else begin
                                                                if (6'h23 == _T_183) begin
                                                                  mem_35 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h23 == _T_178) begin
                                                                    mem_35 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h23 == _T_173) begin
                                                                      mem_35 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h23 == _T_168) begin
                                                                        mem_35 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h23 == _T_163) begin
                                                                          mem_35 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h23 == _T_158) begin
                                                                            mem_35 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h23 == _T_153) begin
                                                                              mem_35 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h23 == _T_308) begin
              mem_35 <= _GEN_31;
            end else begin
              if (6'h23 == _T_303) begin
                mem_35 <= _GEN_30;
              end else begin
                if (6'h23 == _T_298) begin
                  mem_35 <= _GEN_29;
                end else begin
                  if (6'h23 == _T_293) begin
                    mem_35 <= _GEN_28;
                  end else begin
                    if (6'h23 == _T_288) begin
                      mem_35 <= _GEN_27;
                    end else begin
                      if (6'h23 == _T_283) begin
                        mem_35 <= _GEN_26;
                      end else begin
                        if (6'h23 == _T_278) begin
                          mem_35 <= _GEN_25;
                        end else begin
                          if (6'h23 == _T_273) begin
                            mem_35 <= _GEN_24;
                          end else begin
                            if (6'h23 == _T_268) begin
                              mem_35 <= _GEN_23;
                            end else begin
                              if (6'h23 == _T_263) begin
                                mem_35 <= _GEN_22;
                              end else begin
                                if (6'h23 == _T_258) begin
                                  mem_35 <= _GEN_21;
                                end else begin
                                  if (6'h23 == _T_253) begin
                                    mem_35 <= _GEN_20;
                                  end else begin
                                    if (6'h23 == _T_248) begin
                                      mem_35 <= _GEN_19;
                                    end else begin
                                      if (6'h23 == _T_243) begin
                                        mem_35 <= _GEN_18;
                                      end else begin
                                        if (6'h23 == _T_238) begin
                                          mem_35 <= _GEN_17;
                                        end else begin
                                          if (6'h23 == _T_233) begin
                                            mem_35 <= _GEN_16;
                                          end else begin
                                            if (6'h23 == _T_228) begin
                                              mem_35 <= _GEN_15;
                                            end else begin
                                              if (6'h23 == _T_223) begin
                                                mem_35 <= _GEN_14;
                                              end else begin
                                                if (6'h23 == _T_218) begin
                                                  mem_35 <= _GEN_13;
                                                end else begin
                                                  if (6'h23 == _T_213) begin
                                                    mem_35 <= _GEN_12;
                                                  end else begin
                                                    if (6'h23 == _T_208) begin
                                                      mem_35 <= _GEN_11;
                                                    end else begin
                                                      if (6'h23 == _T_203) begin
                                                        mem_35 <= _GEN_10;
                                                      end else begin
                                                        if (6'h23 == _T_198) begin
                                                          mem_35 <= _GEN_9;
                                                        end else begin
                                                          if (6'h23 == _T_193) begin
                                                            mem_35 <= _GEN_8;
                                                          end else begin
                                                            if (6'h23 == _T_188) begin
                                                              mem_35 <= _GEN_7;
                                                            end else begin
                                                              if (6'h23 == _T_183) begin
                                                                mem_35 <= _GEN_6;
                                                              end else begin
                                                                if (6'h23 == _T_178) begin
                                                                  mem_35 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h23 == _T_173) begin
                                                                    mem_35 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h23 == _T_168) begin
                                                                      mem_35 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h23 == _T_163) begin
                                                                        mem_35 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h23 == _T_158) begin
                                                                          mem_35 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h23 == _T_153) begin
                                                                            mem_35 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h23 == _T_308) begin
            mem_35 <= _GEN_31;
          end else begin
            if (6'h23 == _T_303) begin
              mem_35 <= _GEN_30;
            end else begin
              if (6'h23 == _T_298) begin
                mem_35 <= _GEN_29;
              end else begin
                if (6'h23 == _T_293) begin
                  mem_35 <= _GEN_28;
                end else begin
                  if (6'h23 == _T_288) begin
                    mem_35 <= _GEN_27;
                  end else begin
                    if (6'h23 == _T_283) begin
                      mem_35 <= _GEN_26;
                    end else begin
                      if (6'h23 == _T_278) begin
                        mem_35 <= _GEN_25;
                      end else begin
                        if (6'h23 == _T_273) begin
                          mem_35 <= _GEN_24;
                        end else begin
                          if (6'h23 == _T_268) begin
                            mem_35 <= _GEN_23;
                          end else begin
                            if (6'h23 == _T_263) begin
                              mem_35 <= _GEN_22;
                            end else begin
                              if (6'h23 == _T_258) begin
                                mem_35 <= _GEN_21;
                              end else begin
                                if (6'h23 == _T_253) begin
                                  mem_35 <= _GEN_20;
                                end else begin
                                  if (6'h23 == _T_248) begin
                                    mem_35 <= _GEN_19;
                                  end else begin
                                    if (6'h23 == _T_243) begin
                                      mem_35 <= _GEN_18;
                                    end else begin
                                      if (6'h23 == _T_238) begin
                                        mem_35 <= _GEN_17;
                                      end else begin
                                        if (6'h23 == _T_233) begin
                                          mem_35 <= _GEN_16;
                                        end else begin
                                          if (6'h23 == _T_228) begin
                                            mem_35 <= _GEN_15;
                                          end else begin
                                            if (6'h23 == _T_223) begin
                                              mem_35 <= _GEN_14;
                                            end else begin
                                              if (6'h23 == _T_218) begin
                                                mem_35 <= _GEN_13;
                                              end else begin
                                                if (6'h23 == _T_213) begin
                                                  mem_35 <= _GEN_12;
                                                end else begin
                                                  if (6'h23 == _T_208) begin
                                                    mem_35 <= _GEN_11;
                                                  end else begin
                                                    if (6'h23 == _T_203) begin
                                                      mem_35 <= _GEN_10;
                                                    end else begin
                                                      if (6'h23 == _T_198) begin
                                                        mem_35 <= _GEN_9;
                                                      end else begin
                                                        if (6'h23 == _T_193) begin
                                                          mem_35 <= _GEN_8;
                                                        end else begin
                                                          if (6'h23 == _T_188) begin
                                                            mem_35 <= _GEN_7;
                                                          end else begin
                                                            if (6'h23 == _T_183) begin
                                                              mem_35 <= _GEN_6;
                                                            end else begin
                                                              if (6'h23 == _T_178) begin
                                                                mem_35 <= _GEN_5;
                                                              end else begin
                                                                if (6'h23 == _T_173) begin
                                                                  mem_35 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h23 == _T_168) begin
                                                                    mem_35 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h23 == _T_163) begin
                                                                      mem_35 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h23 == _T_158) begin
                                                                        mem_35 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h23 == _T_153) begin
                                                                          mem_35 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h23 == _T_308) begin
          mem_35 <= _GEN_31;
        end else begin
          if (6'h23 == _T_303) begin
            mem_35 <= _GEN_30;
          end else begin
            if (6'h23 == _T_298) begin
              mem_35 <= _GEN_29;
            end else begin
              if (6'h23 == _T_293) begin
                mem_35 <= _GEN_28;
              end else begin
                if (6'h23 == _T_288) begin
                  mem_35 <= _GEN_27;
                end else begin
                  if (6'h23 == _T_283) begin
                    mem_35 <= _GEN_26;
                  end else begin
                    if (6'h23 == _T_278) begin
                      mem_35 <= _GEN_25;
                    end else begin
                      if (6'h23 == _T_273) begin
                        mem_35 <= _GEN_24;
                      end else begin
                        if (6'h23 == _T_268) begin
                          mem_35 <= _GEN_23;
                        end else begin
                          if (6'h23 == _T_263) begin
                            mem_35 <= _GEN_22;
                          end else begin
                            if (6'h23 == _T_258) begin
                              mem_35 <= _GEN_21;
                            end else begin
                              if (6'h23 == _T_253) begin
                                mem_35 <= _GEN_20;
                              end else begin
                                if (6'h23 == _T_248) begin
                                  mem_35 <= _GEN_19;
                                end else begin
                                  if (6'h23 == _T_243) begin
                                    mem_35 <= _GEN_18;
                                  end else begin
                                    if (6'h23 == _T_238) begin
                                      mem_35 <= _GEN_17;
                                    end else begin
                                      if (6'h23 == _T_233) begin
                                        mem_35 <= _GEN_16;
                                      end else begin
                                        if (6'h23 == _T_228) begin
                                          mem_35 <= _GEN_15;
                                        end else begin
                                          if (6'h23 == _T_223) begin
                                            mem_35 <= _GEN_14;
                                          end else begin
                                            if (6'h23 == _T_218) begin
                                              mem_35 <= _GEN_13;
                                            end else begin
                                              if (6'h23 == _T_213) begin
                                                mem_35 <= _GEN_12;
                                              end else begin
                                                if (6'h23 == _T_208) begin
                                                  mem_35 <= _GEN_11;
                                                end else begin
                                                  if (6'h23 == _T_203) begin
                                                    mem_35 <= _GEN_10;
                                                  end else begin
                                                    if (6'h23 == _T_198) begin
                                                      mem_35 <= _GEN_9;
                                                    end else begin
                                                      if (6'h23 == _T_193) begin
                                                        mem_35 <= _GEN_8;
                                                      end else begin
                                                        if (6'h23 == _T_188) begin
                                                          mem_35 <= _GEN_7;
                                                        end else begin
                                                          if (6'h23 == _T_183) begin
                                                            mem_35 <= _GEN_6;
                                                          end else begin
                                                            if (6'h23 == _T_178) begin
                                                              mem_35 <= _GEN_5;
                                                            end else begin
                                                              if (6'h23 == _T_173) begin
                                                                mem_35 <= _GEN_4;
                                                              end else begin
                                                                if (6'h23 == _T_168) begin
                                                                  mem_35 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h23 == _T_163) begin
                                                                    mem_35 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h23 == _T_158) begin
                                                                      mem_35 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h23 == _T_153) begin
                                                                        mem_35 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h24 == wPos) begin
            mem_36 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h24 == _T_308) begin
                mem_36 <= _GEN_31;
              end else begin
                if (6'h24 == _T_303) begin
                  mem_36 <= _GEN_30;
                end else begin
                  if (6'h24 == _T_298) begin
                    mem_36 <= _GEN_29;
                  end else begin
                    if (6'h24 == _T_293) begin
                      mem_36 <= _GEN_28;
                    end else begin
                      if (6'h24 == _T_288) begin
                        mem_36 <= _GEN_27;
                      end else begin
                        if (6'h24 == _T_283) begin
                          mem_36 <= _GEN_26;
                        end else begin
                          if (6'h24 == _T_278) begin
                            mem_36 <= _GEN_25;
                          end else begin
                            if (6'h24 == _T_273) begin
                              mem_36 <= _GEN_24;
                            end else begin
                              if (6'h24 == _T_268) begin
                                mem_36 <= _GEN_23;
                              end else begin
                                if (6'h24 == _T_263) begin
                                  mem_36 <= _GEN_22;
                                end else begin
                                  if (6'h24 == _T_258) begin
                                    mem_36 <= _GEN_21;
                                  end else begin
                                    if (6'h24 == _T_253) begin
                                      mem_36 <= _GEN_20;
                                    end else begin
                                      if (6'h24 == _T_248) begin
                                        mem_36 <= _GEN_19;
                                      end else begin
                                        if (6'h24 == _T_243) begin
                                          mem_36 <= _GEN_18;
                                        end else begin
                                          if (6'h24 == _T_238) begin
                                            mem_36 <= _GEN_17;
                                          end else begin
                                            if (6'h24 == _T_233) begin
                                              mem_36 <= _GEN_16;
                                            end else begin
                                              if (6'h24 == _T_228) begin
                                                mem_36 <= _GEN_15;
                                              end else begin
                                                if (6'h24 == _T_223) begin
                                                  mem_36 <= _GEN_14;
                                                end else begin
                                                  if (6'h24 == _T_218) begin
                                                    mem_36 <= _GEN_13;
                                                  end else begin
                                                    if (6'h24 == _T_213) begin
                                                      mem_36 <= _GEN_12;
                                                    end else begin
                                                      if (6'h24 == _T_208) begin
                                                        mem_36 <= _GEN_11;
                                                      end else begin
                                                        if (6'h24 == _T_203) begin
                                                          mem_36 <= _GEN_10;
                                                        end else begin
                                                          if (6'h24 == _T_198) begin
                                                            mem_36 <= _GEN_9;
                                                          end else begin
                                                            if (6'h24 == _T_193) begin
                                                              mem_36 <= _GEN_8;
                                                            end else begin
                                                              if (6'h24 == _T_188) begin
                                                                mem_36 <= _GEN_7;
                                                              end else begin
                                                                if (6'h24 == _T_183) begin
                                                                  mem_36 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h24 == _T_178) begin
                                                                    mem_36 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h24 == _T_173) begin
                                                                      mem_36 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h24 == _T_168) begin
                                                                        mem_36 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h24 == _T_163) begin
                                                                          mem_36 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h24 == _T_158) begin
                                                                            mem_36 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h24 == _T_153) begin
                                                                              mem_36 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h24 == _T_308) begin
              mem_36 <= _GEN_31;
            end else begin
              if (6'h24 == _T_303) begin
                mem_36 <= _GEN_30;
              end else begin
                if (6'h24 == _T_298) begin
                  mem_36 <= _GEN_29;
                end else begin
                  if (6'h24 == _T_293) begin
                    mem_36 <= _GEN_28;
                  end else begin
                    if (6'h24 == _T_288) begin
                      mem_36 <= _GEN_27;
                    end else begin
                      if (6'h24 == _T_283) begin
                        mem_36 <= _GEN_26;
                      end else begin
                        if (6'h24 == _T_278) begin
                          mem_36 <= _GEN_25;
                        end else begin
                          if (6'h24 == _T_273) begin
                            mem_36 <= _GEN_24;
                          end else begin
                            if (6'h24 == _T_268) begin
                              mem_36 <= _GEN_23;
                            end else begin
                              if (6'h24 == _T_263) begin
                                mem_36 <= _GEN_22;
                              end else begin
                                if (6'h24 == _T_258) begin
                                  mem_36 <= _GEN_21;
                                end else begin
                                  if (6'h24 == _T_253) begin
                                    mem_36 <= _GEN_20;
                                  end else begin
                                    if (6'h24 == _T_248) begin
                                      mem_36 <= _GEN_19;
                                    end else begin
                                      if (6'h24 == _T_243) begin
                                        mem_36 <= _GEN_18;
                                      end else begin
                                        if (6'h24 == _T_238) begin
                                          mem_36 <= _GEN_17;
                                        end else begin
                                          if (6'h24 == _T_233) begin
                                            mem_36 <= _GEN_16;
                                          end else begin
                                            if (6'h24 == _T_228) begin
                                              mem_36 <= _GEN_15;
                                            end else begin
                                              if (6'h24 == _T_223) begin
                                                mem_36 <= _GEN_14;
                                              end else begin
                                                if (6'h24 == _T_218) begin
                                                  mem_36 <= _GEN_13;
                                                end else begin
                                                  if (6'h24 == _T_213) begin
                                                    mem_36 <= _GEN_12;
                                                  end else begin
                                                    if (6'h24 == _T_208) begin
                                                      mem_36 <= _GEN_11;
                                                    end else begin
                                                      if (6'h24 == _T_203) begin
                                                        mem_36 <= _GEN_10;
                                                      end else begin
                                                        if (6'h24 == _T_198) begin
                                                          mem_36 <= _GEN_9;
                                                        end else begin
                                                          if (6'h24 == _T_193) begin
                                                            mem_36 <= _GEN_8;
                                                          end else begin
                                                            if (6'h24 == _T_188) begin
                                                              mem_36 <= _GEN_7;
                                                            end else begin
                                                              if (6'h24 == _T_183) begin
                                                                mem_36 <= _GEN_6;
                                                              end else begin
                                                                if (6'h24 == _T_178) begin
                                                                  mem_36 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h24 == _T_173) begin
                                                                    mem_36 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h24 == _T_168) begin
                                                                      mem_36 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h24 == _T_163) begin
                                                                        mem_36 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h24 == _T_158) begin
                                                                          mem_36 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h24 == _T_153) begin
                                                                            mem_36 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h24 == _T_308) begin
            mem_36 <= _GEN_31;
          end else begin
            if (6'h24 == _T_303) begin
              mem_36 <= _GEN_30;
            end else begin
              if (6'h24 == _T_298) begin
                mem_36 <= _GEN_29;
              end else begin
                if (6'h24 == _T_293) begin
                  mem_36 <= _GEN_28;
                end else begin
                  if (6'h24 == _T_288) begin
                    mem_36 <= _GEN_27;
                  end else begin
                    if (6'h24 == _T_283) begin
                      mem_36 <= _GEN_26;
                    end else begin
                      if (6'h24 == _T_278) begin
                        mem_36 <= _GEN_25;
                      end else begin
                        if (6'h24 == _T_273) begin
                          mem_36 <= _GEN_24;
                        end else begin
                          if (6'h24 == _T_268) begin
                            mem_36 <= _GEN_23;
                          end else begin
                            if (6'h24 == _T_263) begin
                              mem_36 <= _GEN_22;
                            end else begin
                              if (6'h24 == _T_258) begin
                                mem_36 <= _GEN_21;
                              end else begin
                                if (6'h24 == _T_253) begin
                                  mem_36 <= _GEN_20;
                                end else begin
                                  if (6'h24 == _T_248) begin
                                    mem_36 <= _GEN_19;
                                  end else begin
                                    if (6'h24 == _T_243) begin
                                      mem_36 <= _GEN_18;
                                    end else begin
                                      if (6'h24 == _T_238) begin
                                        mem_36 <= _GEN_17;
                                      end else begin
                                        if (6'h24 == _T_233) begin
                                          mem_36 <= _GEN_16;
                                        end else begin
                                          if (6'h24 == _T_228) begin
                                            mem_36 <= _GEN_15;
                                          end else begin
                                            if (6'h24 == _T_223) begin
                                              mem_36 <= _GEN_14;
                                            end else begin
                                              if (6'h24 == _T_218) begin
                                                mem_36 <= _GEN_13;
                                              end else begin
                                                if (6'h24 == _T_213) begin
                                                  mem_36 <= _GEN_12;
                                                end else begin
                                                  if (6'h24 == _T_208) begin
                                                    mem_36 <= _GEN_11;
                                                  end else begin
                                                    if (6'h24 == _T_203) begin
                                                      mem_36 <= _GEN_10;
                                                    end else begin
                                                      if (6'h24 == _T_198) begin
                                                        mem_36 <= _GEN_9;
                                                      end else begin
                                                        if (6'h24 == _T_193) begin
                                                          mem_36 <= _GEN_8;
                                                        end else begin
                                                          if (6'h24 == _T_188) begin
                                                            mem_36 <= _GEN_7;
                                                          end else begin
                                                            if (6'h24 == _T_183) begin
                                                              mem_36 <= _GEN_6;
                                                            end else begin
                                                              if (6'h24 == _T_178) begin
                                                                mem_36 <= _GEN_5;
                                                              end else begin
                                                                if (6'h24 == _T_173) begin
                                                                  mem_36 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h24 == _T_168) begin
                                                                    mem_36 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h24 == _T_163) begin
                                                                      mem_36 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h24 == _T_158) begin
                                                                        mem_36 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h24 == _T_153) begin
                                                                          mem_36 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h24 == _T_308) begin
          mem_36 <= _GEN_31;
        end else begin
          if (6'h24 == _T_303) begin
            mem_36 <= _GEN_30;
          end else begin
            if (6'h24 == _T_298) begin
              mem_36 <= _GEN_29;
            end else begin
              if (6'h24 == _T_293) begin
                mem_36 <= _GEN_28;
              end else begin
                if (6'h24 == _T_288) begin
                  mem_36 <= _GEN_27;
                end else begin
                  if (6'h24 == _T_283) begin
                    mem_36 <= _GEN_26;
                  end else begin
                    if (6'h24 == _T_278) begin
                      mem_36 <= _GEN_25;
                    end else begin
                      if (6'h24 == _T_273) begin
                        mem_36 <= _GEN_24;
                      end else begin
                        if (6'h24 == _T_268) begin
                          mem_36 <= _GEN_23;
                        end else begin
                          if (6'h24 == _T_263) begin
                            mem_36 <= _GEN_22;
                          end else begin
                            if (6'h24 == _T_258) begin
                              mem_36 <= _GEN_21;
                            end else begin
                              if (6'h24 == _T_253) begin
                                mem_36 <= _GEN_20;
                              end else begin
                                if (6'h24 == _T_248) begin
                                  mem_36 <= _GEN_19;
                                end else begin
                                  if (6'h24 == _T_243) begin
                                    mem_36 <= _GEN_18;
                                  end else begin
                                    if (6'h24 == _T_238) begin
                                      mem_36 <= _GEN_17;
                                    end else begin
                                      if (6'h24 == _T_233) begin
                                        mem_36 <= _GEN_16;
                                      end else begin
                                        if (6'h24 == _T_228) begin
                                          mem_36 <= _GEN_15;
                                        end else begin
                                          if (6'h24 == _T_223) begin
                                            mem_36 <= _GEN_14;
                                          end else begin
                                            if (6'h24 == _T_218) begin
                                              mem_36 <= _GEN_13;
                                            end else begin
                                              if (6'h24 == _T_213) begin
                                                mem_36 <= _GEN_12;
                                              end else begin
                                                if (6'h24 == _T_208) begin
                                                  mem_36 <= _GEN_11;
                                                end else begin
                                                  if (6'h24 == _T_203) begin
                                                    mem_36 <= _GEN_10;
                                                  end else begin
                                                    if (6'h24 == _T_198) begin
                                                      mem_36 <= _GEN_9;
                                                    end else begin
                                                      if (6'h24 == _T_193) begin
                                                        mem_36 <= _GEN_8;
                                                      end else begin
                                                        if (6'h24 == _T_188) begin
                                                          mem_36 <= _GEN_7;
                                                        end else begin
                                                          if (6'h24 == _T_183) begin
                                                            mem_36 <= _GEN_6;
                                                          end else begin
                                                            if (6'h24 == _T_178) begin
                                                              mem_36 <= _GEN_5;
                                                            end else begin
                                                              if (6'h24 == _T_173) begin
                                                                mem_36 <= _GEN_4;
                                                              end else begin
                                                                if (6'h24 == _T_168) begin
                                                                  mem_36 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h24 == _T_163) begin
                                                                    mem_36 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h24 == _T_158) begin
                                                                      mem_36 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h24 == _T_153) begin
                                                                        mem_36 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h25 == wPos) begin
            mem_37 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h25 == _T_308) begin
                mem_37 <= _GEN_31;
              end else begin
                if (6'h25 == _T_303) begin
                  mem_37 <= _GEN_30;
                end else begin
                  if (6'h25 == _T_298) begin
                    mem_37 <= _GEN_29;
                  end else begin
                    if (6'h25 == _T_293) begin
                      mem_37 <= _GEN_28;
                    end else begin
                      if (6'h25 == _T_288) begin
                        mem_37 <= _GEN_27;
                      end else begin
                        if (6'h25 == _T_283) begin
                          mem_37 <= _GEN_26;
                        end else begin
                          if (6'h25 == _T_278) begin
                            mem_37 <= _GEN_25;
                          end else begin
                            if (6'h25 == _T_273) begin
                              mem_37 <= _GEN_24;
                            end else begin
                              if (6'h25 == _T_268) begin
                                mem_37 <= _GEN_23;
                              end else begin
                                if (6'h25 == _T_263) begin
                                  mem_37 <= _GEN_22;
                                end else begin
                                  if (6'h25 == _T_258) begin
                                    mem_37 <= _GEN_21;
                                  end else begin
                                    if (6'h25 == _T_253) begin
                                      mem_37 <= _GEN_20;
                                    end else begin
                                      if (6'h25 == _T_248) begin
                                        mem_37 <= _GEN_19;
                                      end else begin
                                        if (6'h25 == _T_243) begin
                                          mem_37 <= _GEN_18;
                                        end else begin
                                          if (6'h25 == _T_238) begin
                                            mem_37 <= _GEN_17;
                                          end else begin
                                            if (6'h25 == _T_233) begin
                                              mem_37 <= _GEN_16;
                                            end else begin
                                              if (6'h25 == _T_228) begin
                                                mem_37 <= _GEN_15;
                                              end else begin
                                                if (6'h25 == _T_223) begin
                                                  mem_37 <= _GEN_14;
                                                end else begin
                                                  if (6'h25 == _T_218) begin
                                                    mem_37 <= _GEN_13;
                                                  end else begin
                                                    if (6'h25 == _T_213) begin
                                                      mem_37 <= _GEN_12;
                                                    end else begin
                                                      if (6'h25 == _T_208) begin
                                                        mem_37 <= _GEN_11;
                                                      end else begin
                                                        if (6'h25 == _T_203) begin
                                                          mem_37 <= _GEN_10;
                                                        end else begin
                                                          if (6'h25 == _T_198) begin
                                                            mem_37 <= _GEN_9;
                                                          end else begin
                                                            if (6'h25 == _T_193) begin
                                                              mem_37 <= _GEN_8;
                                                            end else begin
                                                              if (6'h25 == _T_188) begin
                                                                mem_37 <= _GEN_7;
                                                              end else begin
                                                                if (6'h25 == _T_183) begin
                                                                  mem_37 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h25 == _T_178) begin
                                                                    mem_37 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h25 == _T_173) begin
                                                                      mem_37 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h25 == _T_168) begin
                                                                        mem_37 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h25 == _T_163) begin
                                                                          mem_37 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h25 == _T_158) begin
                                                                            mem_37 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h25 == _T_153) begin
                                                                              mem_37 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h25 == _T_308) begin
              mem_37 <= _GEN_31;
            end else begin
              if (6'h25 == _T_303) begin
                mem_37 <= _GEN_30;
              end else begin
                if (6'h25 == _T_298) begin
                  mem_37 <= _GEN_29;
                end else begin
                  if (6'h25 == _T_293) begin
                    mem_37 <= _GEN_28;
                  end else begin
                    if (6'h25 == _T_288) begin
                      mem_37 <= _GEN_27;
                    end else begin
                      if (6'h25 == _T_283) begin
                        mem_37 <= _GEN_26;
                      end else begin
                        if (6'h25 == _T_278) begin
                          mem_37 <= _GEN_25;
                        end else begin
                          if (6'h25 == _T_273) begin
                            mem_37 <= _GEN_24;
                          end else begin
                            if (6'h25 == _T_268) begin
                              mem_37 <= _GEN_23;
                            end else begin
                              if (6'h25 == _T_263) begin
                                mem_37 <= _GEN_22;
                              end else begin
                                if (6'h25 == _T_258) begin
                                  mem_37 <= _GEN_21;
                                end else begin
                                  if (6'h25 == _T_253) begin
                                    mem_37 <= _GEN_20;
                                  end else begin
                                    if (6'h25 == _T_248) begin
                                      mem_37 <= _GEN_19;
                                    end else begin
                                      if (6'h25 == _T_243) begin
                                        mem_37 <= _GEN_18;
                                      end else begin
                                        if (6'h25 == _T_238) begin
                                          mem_37 <= _GEN_17;
                                        end else begin
                                          if (6'h25 == _T_233) begin
                                            mem_37 <= _GEN_16;
                                          end else begin
                                            if (6'h25 == _T_228) begin
                                              mem_37 <= _GEN_15;
                                            end else begin
                                              if (6'h25 == _T_223) begin
                                                mem_37 <= _GEN_14;
                                              end else begin
                                                if (6'h25 == _T_218) begin
                                                  mem_37 <= _GEN_13;
                                                end else begin
                                                  if (6'h25 == _T_213) begin
                                                    mem_37 <= _GEN_12;
                                                  end else begin
                                                    if (6'h25 == _T_208) begin
                                                      mem_37 <= _GEN_11;
                                                    end else begin
                                                      if (6'h25 == _T_203) begin
                                                        mem_37 <= _GEN_10;
                                                      end else begin
                                                        if (6'h25 == _T_198) begin
                                                          mem_37 <= _GEN_9;
                                                        end else begin
                                                          if (6'h25 == _T_193) begin
                                                            mem_37 <= _GEN_8;
                                                          end else begin
                                                            if (6'h25 == _T_188) begin
                                                              mem_37 <= _GEN_7;
                                                            end else begin
                                                              if (6'h25 == _T_183) begin
                                                                mem_37 <= _GEN_6;
                                                              end else begin
                                                                if (6'h25 == _T_178) begin
                                                                  mem_37 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h25 == _T_173) begin
                                                                    mem_37 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h25 == _T_168) begin
                                                                      mem_37 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h25 == _T_163) begin
                                                                        mem_37 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h25 == _T_158) begin
                                                                          mem_37 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h25 == _T_153) begin
                                                                            mem_37 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h25 == _T_308) begin
            mem_37 <= _GEN_31;
          end else begin
            if (6'h25 == _T_303) begin
              mem_37 <= _GEN_30;
            end else begin
              if (6'h25 == _T_298) begin
                mem_37 <= _GEN_29;
              end else begin
                if (6'h25 == _T_293) begin
                  mem_37 <= _GEN_28;
                end else begin
                  if (6'h25 == _T_288) begin
                    mem_37 <= _GEN_27;
                  end else begin
                    if (6'h25 == _T_283) begin
                      mem_37 <= _GEN_26;
                    end else begin
                      if (6'h25 == _T_278) begin
                        mem_37 <= _GEN_25;
                      end else begin
                        if (6'h25 == _T_273) begin
                          mem_37 <= _GEN_24;
                        end else begin
                          if (6'h25 == _T_268) begin
                            mem_37 <= _GEN_23;
                          end else begin
                            if (6'h25 == _T_263) begin
                              mem_37 <= _GEN_22;
                            end else begin
                              if (6'h25 == _T_258) begin
                                mem_37 <= _GEN_21;
                              end else begin
                                if (6'h25 == _T_253) begin
                                  mem_37 <= _GEN_20;
                                end else begin
                                  if (6'h25 == _T_248) begin
                                    mem_37 <= _GEN_19;
                                  end else begin
                                    if (6'h25 == _T_243) begin
                                      mem_37 <= _GEN_18;
                                    end else begin
                                      if (6'h25 == _T_238) begin
                                        mem_37 <= _GEN_17;
                                      end else begin
                                        if (6'h25 == _T_233) begin
                                          mem_37 <= _GEN_16;
                                        end else begin
                                          if (6'h25 == _T_228) begin
                                            mem_37 <= _GEN_15;
                                          end else begin
                                            if (6'h25 == _T_223) begin
                                              mem_37 <= _GEN_14;
                                            end else begin
                                              if (6'h25 == _T_218) begin
                                                mem_37 <= _GEN_13;
                                              end else begin
                                                if (6'h25 == _T_213) begin
                                                  mem_37 <= _GEN_12;
                                                end else begin
                                                  if (6'h25 == _T_208) begin
                                                    mem_37 <= _GEN_11;
                                                  end else begin
                                                    if (6'h25 == _T_203) begin
                                                      mem_37 <= _GEN_10;
                                                    end else begin
                                                      if (6'h25 == _T_198) begin
                                                        mem_37 <= _GEN_9;
                                                      end else begin
                                                        if (6'h25 == _T_193) begin
                                                          mem_37 <= _GEN_8;
                                                        end else begin
                                                          if (6'h25 == _T_188) begin
                                                            mem_37 <= _GEN_7;
                                                          end else begin
                                                            if (6'h25 == _T_183) begin
                                                              mem_37 <= _GEN_6;
                                                            end else begin
                                                              if (6'h25 == _T_178) begin
                                                                mem_37 <= _GEN_5;
                                                              end else begin
                                                                if (6'h25 == _T_173) begin
                                                                  mem_37 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h25 == _T_168) begin
                                                                    mem_37 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h25 == _T_163) begin
                                                                      mem_37 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h25 == _T_158) begin
                                                                        mem_37 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h25 == _T_153) begin
                                                                          mem_37 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h25 == _T_308) begin
          mem_37 <= _GEN_31;
        end else begin
          if (6'h25 == _T_303) begin
            mem_37 <= _GEN_30;
          end else begin
            if (6'h25 == _T_298) begin
              mem_37 <= _GEN_29;
            end else begin
              if (6'h25 == _T_293) begin
                mem_37 <= _GEN_28;
              end else begin
                if (6'h25 == _T_288) begin
                  mem_37 <= _GEN_27;
                end else begin
                  if (6'h25 == _T_283) begin
                    mem_37 <= _GEN_26;
                  end else begin
                    if (6'h25 == _T_278) begin
                      mem_37 <= _GEN_25;
                    end else begin
                      if (6'h25 == _T_273) begin
                        mem_37 <= _GEN_24;
                      end else begin
                        if (6'h25 == _T_268) begin
                          mem_37 <= _GEN_23;
                        end else begin
                          if (6'h25 == _T_263) begin
                            mem_37 <= _GEN_22;
                          end else begin
                            if (6'h25 == _T_258) begin
                              mem_37 <= _GEN_21;
                            end else begin
                              if (6'h25 == _T_253) begin
                                mem_37 <= _GEN_20;
                              end else begin
                                if (6'h25 == _T_248) begin
                                  mem_37 <= _GEN_19;
                                end else begin
                                  if (6'h25 == _T_243) begin
                                    mem_37 <= _GEN_18;
                                  end else begin
                                    if (6'h25 == _T_238) begin
                                      mem_37 <= _GEN_17;
                                    end else begin
                                      if (6'h25 == _T_233) begin
                                        mem_37 <= _GEN_16;
                                      end else begin
                                        if (6'h25 == _T_228) begin
                                          mem_37 <= _GEN_15;
                                        end else begin
                                          if (6'h25 == _T_223) begin
                                            mem_37 <= _GEN_14;
                                          end else begin
                                            if (6'h25 == _T_218) begin
                                              mem_37 <= _GEN_13;
                                            end else begin
                                              if (6'h25 == _T_213) begin
                                                mem_37 <= _GEN_12;
                                              end else begin
                                                if (6'h25 == _T_208) begin
                                                  mem_37 <= _GEN_11;
                                                end else begin
                                                  if (6'h25 == _T_203) begin
                                                    mem_37 <= _GEN_10;
                                                  end else begin
                                                    if (6'h25 == _T_198) begin
                                                      mem_37 <= _GEN_9;
                                                    end else begin
                                                      if (6'h25 == _T_193) begin
                                                        mem_37 <= _GEN_8;
                                                      end else begin
                                                        if (6'h25 == _T_188) begin
                                                          mem_37 <= _GEN_7;
                                                        end else begin
                                                          if (6'h25 == _T_183) begin
                                                            mem_37 <= _GEN_6;
                                                          end else begin
                                                            if (6'h25 == _T_178) begin
                                                              mem_37 <= _GEN_5;
                                                            end else begin
                                                              if (6'h25 == _T_173) begin
                                                                mem_37 <= _GEN_4;
                                                              end else begin
                                                                if (6'h25 == _T_168) begin
                                                                  mem_37 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h25 == _T_163) begin
                                                                    mem_37 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h25 == _T_158) begin
                                                                      mem_37 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h25 == _T_153) begin
                                                                        mem_37 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h26 == wPos) begin
            mem_38 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h26 == _T_308) begin
                mem_38 <= _GEN_31;
              end else begin
                if (6'h26 == _T_303) begin
                  mem_38 <= _GEN_30;
                end else begin
                  if (6'h26 == _T_298) begin
                    mem_38 <= _GEN_29;
                  end else begin
                    if (6'h26 == _T_293) begin
                      mem_38 <= _GEN_28;
                    end else begin
                      if (6'h26 == _T_288) begin
                        mem_38 <= _GEN_27;
                      end else begin
                        if (6'h26 == _T_283) begin
                          mem_38 <= _GEN_26;
                        end else begin
                          if (6'h26 == _T_278) begin
                            mem_38 <= _GEN_25;
                          end else begin
                            if (6'h26 == _T_273) begin
                              mem_38 <= _GEN_24;
                            end else begin
                              if (6'h26 == _T_268) begin
                                mem_38 <= _GEN_23;
                              end else begin
                                if (6'h26 == _T_263) begin
                                  mem_38 <= _GEN_22;
                                end else begin
                                  if (6'h26 == _T_258) begin
                                    mem_38 <= _GEN_21;
                                  end else begin
                                    if (6'h26 == _T_253) begin
                                      mem_38 <= _GEN_20;
                                    end else begin
                                      if (6'h26 == _T_248) begin
                                        mem_38 <= _GEN_19;
                                      end else begin
                                        if (6'h26 == _T_243) begin
                                          mem_38 <= _GEN_18;
                                        end else begin
                                          if (6'h26 == _T_238) begin
                                            mem_38 <= _GEN_17;
                                          end else begin
                                            if (6'h26 == _T_233) begin
                                              mem_38 <= _GEN_16;
                                            end else begin
                                              if (6'h26 == _T_228) begin
                                                mem_38 <= _GEN_15;
                                              end else begin
                                                if (6'h26 == _T_223) begin
                                                  mem_38 <= _GEN_14;
                                                end else begin
                                                  if (6'h26 == _T_218) begin
                                                    mem_38 <= _GEN_13;
                                                  end else begin
                                                    if (6'h26 == _T_213) begin
                                                      mem_38 <= _GEN_12;
                                                    end else begin
                                                      if (6'h26 == _T_208) begin
                                                        mem_38 <= _GEN_11;
                                                      end else begin
                                                        if (6'h26 == _T_203) begin
                                                          mem_38 <= _GEN_10;
                                                        end else begin
                                                          if (6'h26 == _T_198) begin
                                                            mem_38 <= _GEN_9;
                                                          end else begin
                                                            if (6'h26 == _T_193) begin
                                                              mem_38 <= _GEN_8;
                                                            end else begin
                                                              if (6'h26 == _T_188) begin
                                                                mem_38 <= _GEN_7;
                                                              end else begin
                                                                if (6'h26 == _T_183) begin
                                                                  mem_38 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h26 == _T_178) begin
                                                                    mem_38 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h26 == _T_173) begin
                                                                      mem_38 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h26 == _T_168) begin
                                                                        mem_38 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h26 == _T_163) begin
                                                                          mem_38 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h26 == _T_158) begin
                                                                            mem_38 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h26 == _T_153) begin
                                                                              mem_38 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h26 == _T_308) begin
              mem_38 <= _GEN_31;
            end else begin
              if (6'h26 == _T_303) begin
                mem_38 <= _GEN_30;
              end else begin
                if (6'h26 == _T_298) begin
                  mem_38 <= _GEN_29;
                end else begin
                  if (6'h26 == _T_293) begin
                    mem_38 <= _GEN_28;
                  end else begin
                    if (6'h26 == _T_288) begin
                      mem_38 <= _GEN_27;
                    end else begin
                      if (6'h26 == _T_283) begin
                        mem_38 <= _GEN_26;
                      end else begin
                        if (6'h26 == _T_278) begin
                          mem_38 <= _GEN_25;
                        end else begin
                          if (6'h26 == _T_273) begin
                            mem_38 <= _GEN_24;
                          end else begin
                            if (6'h26 == _T_268) begin
                              mem_38 <= _GEN_23;
                            end else begin
                              if (6'h26 == _T_263) begin
                                mem_38 <= _GEN_22;
                              end else begin
                                if (6'h26 == _T_258) begin
                                  mem_38 <= _GEN_21;
                                end else begin
                                  if (6'h26 == _T_253) begin
                                    mem_38 <= _GEN_20;
                                  end else begin
                                    if (6'h26 == _T_248) begin
                                      mem_38 <= _GEN_19;
                                    end else begin
                                      if (6'h26 == _T_243) begin
                                        mem_38 <= _GEN_18;
                                      end else begin
                                        if (6'h26 == _T_238) begin
                                          mem_38 <= _GEN_17;
                                        end else begin
                                          if (6'h26 == _T_233) begin
                                            mem_38 <= _GEN_16;
                                          end else begin
                                            if (6'h26 == _T_228) begin
                                              mem_38 <= _GEN_15;
                                            end else begin
                                              if (6'h26 == _T_223) begin
                                                mem_38 <= _GEN_14;
                                              end else begin
                                                if (6'h26 == _T_218) begin
                                                  mem_38 <= _GEN_13;
                                                end else begin
                                                  if (6'h26 == _T_213) begin
                                                    mem_38 <= _GEN_12;
                                                  end else begin
                                                    if (6'h26 == _T_208) begin
                                                      mem_38 <= _GEN_11;
                                                    end else begin
                                                      if (6'h26 == _T_203) begin
                                                        mem_38 <= _GEN_10;
                                                      end else begin
                                                        if (6'h26 == _T_198) begin
                                                          mem_38 <= _GEN_9;
                                                        end else begin
                                                          if (6'h26 == _T_193) begin
                                                            mem_38 <= _GEN_8;
                                                          end else begin
                                                            if (6'h26 == _T_188) begin
                                                              mem_38 <= _GEN_7;
                                                            end else begin
                                                              if (6'h26 == _T_183) begin
                                                                mem_38 <= _GEN_6;
                                                              end else begin
                                                                if (6'h26 == _T_178) begin
                                                                  mem_38 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h26 == _T_173) begin
                                                                    mem_38 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h26 == _T_168) begin
                                                                      mem_38 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h26 == _T_163) begin
                                                                        mem_38 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h26 == _T_158) begin
                                                                          mem_38 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h26 == _T_153) begin
                                                                            mem_38 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h26 == _T_308) begin
            mem_38 <= _GEN_31;
          end else begin
            if (6'h26 == _T_303) begin
              mem_38 <= _GEN_30;
            end else begin
              if (6'h26 == _T_298) begin
                mem_38 <= _GEN_29;
              end else begin
                if (6'h26 == _T_293) begin
                  mem_38 <= _GEN_28;
                end else begin
                  if (6'h26 == _T_288) begin
                    mem_38 <= _GEN_27;
                  end else begin
                    if (6'h26 == _T_283) begin
                      mem_38 <= _GEN_26;
                    end else begin
                      if (6'h26 == _T_278) begin
                        mem_38 <= _GEN_25;
                      end else begin
                        if (6'h26 == _T_273) begin
                          mem_38 <= _GEN_24;
                        end else begin
                          if (6'h26 == _T_268) begin
                            mem_38 <= _GEN_23;
                          end else begin
                            if (6'h26 == _T_263) begin
                              mem_38 <= _GEN_22;
                            end else begin
                              if (6'h26 == _T_258) begin
                                mem_38 <= _GEN_21;
                              end else begin
                                if (6'h26 == _T_253) begin
                                  mem_38 <= _GEN_20;
                                end else begin
                                  if (6'h26 == _T_248) begin
                                    mem_38 <= _GEN_19;
                                  end else begin
                                    if (6'h26 == _T_243) begin
                                      mem_38 <= _GEN_18;
                                    end else begin
                                      if (6'h26 == _T_238) begin
                                        mem_38 <= _GEN_17;
                                      end else begin
                                        if (6'h26 == _T_233) begin
                                          mem_38 <= _GEN_16;
                                        end else begin
                                          if (6'h26 == _T_228) begin
                                            mem_38 <= _GEN_15;
                                          end else begin
                                            if (6'h26 == _T_223) begin
                                              mem_38 <= _GEN_14;
                                            end else begin
                                              if (6'h26 == _T_218) begin
                                                mem_38 <= _GEN_13;
                                              end else begin
                                                if (6'h26 == _T_213) begin
                                                  mem_38 <= _GEN_12;
                                                end else begin
                                                  if (6'h26 == _T_208) begin
                                                    mem_38 <= _GEN_11;
                                                  end else begin
                                                    if (6'h26 == _T_203) begin
                                                      mem_38 <= _GEN_10;
                                                    end else begin
                                                      if (6'h26 == _T_198) begin
                                                        mem_38 <= _GEN_9;
                                                      end else begin
                                                        if (6'h26 == _T_193) begin
                                                          mem_38 <= _GEN_8;
                                                        end else begin
                                                          if (6'h26 == _T_188) begin
                                                            mem_38 <= _GEN_7;
                                                          end else begin
                                                            if (6'h26 == _T_183) begin
                                                              mem_38 <= _GEN_6;
                                                            end else begin
                                                              if (6'h26 == _T_178) begin
                                                                mem_38 <= _GEN_5;
                                                              end else begin
                                                                if (6'h26 == _T_173) begin
                                                                  mem_38 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h26 == _T_168) begin
                                                                    mem_38 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h26 == _T_163) begin
                                                                      mem_38 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h26 == _T_158) begin
                                                                        mem_38 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h26 == _T_153) begin
                                                                          mem_38 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h26 == _T_308) begin
          mem_38 <= _GEN_31;
        end else begin
          if (6'h26 == _T_303) begin
            mem_38 <= _GEN_30;
          end else begin
            if (6'h26 == _T_298) begin
              mem_38 <= _GEN_29;
            end else begin
              if (6'h26 == _T_293) begin
                mem_38 <= _GEN_28;
              end else begin
                if (6'h26 == _T_288) begin
                  mem_38 <= _GEN_27;
                end else begin
                  if (6'h26 == _T_283) begin
                    mem_38 <= _GEN_26;
                  end else begin
                    if (6'h26 == _T_278) begin
                      mem_38 <= _GEN_25;
                    end else begin
                      if (6'h26 == _T_273) begin
                        mem_38 <= _GEN_24;
                      end else begin
                        if (6'h26 == _T_268) begin
                          mem_38 <= _GEN_23;
                        end else begin
                          if (6'h26 == _T_263) begin
                            mem_38 <= _GEN_22;
                          end else begin
                            if (6'h26 == _T_258) begin
                              mem_38 <= _GEN_21;
                            end else begin
                              if (6'h26 == _T_253) begin
                                mem_38 <= _GEN_20;
                              end else begin
                                if (6'h26 == _T_248) begin
                                  mem_38 <= _GEN_19;
                                end else begin
                                  if (6'h26 == _T_243) begin
                                    mem_38 <= _GEN_18;
                                  end else begin
                                    if (6'h26 == _T_238) begin
                                      mem_38 <= _GEN_17;
                                    end else begin
                                      if (6'h26 == _T_233) begin
                                        mem_38 <= _GEN_16;
                                      end else begin
                                        if (6'h26 == _T_228) begin
                                          mem_38 <= _GEN_15;
                                        end else begin
                                          if (6'h26 == _T_223) begin
                                            mem_38 <= _GEN_14;
                                          end else begin
                                            if (6'h26 == _T_218) begin
                                              mem_38 <= _GEN_13;
                                            end else begin
                                              if (6'h26 == _T_213) begin
                                                mem_38 <= _GEN_12;
                                              end else begin
                                                if (6'h26 == _T_208) begin
                                                  mem_38 <= _GEN_11;
                                                end else begin
                                                  if (6'h26 == _T_203) begin
                                                    mem_38 <= _GEN_10;
                                                  end else begin
                                                    if (6'h26 == _T_198) begin
                                                      mem_38 <= _GEN_9;
                                                    end else begin
                                                      if (6'h26 == _T_193) begin
                                                        mem_38 <= _GEN_8;
                                                      end else begin
                                                        if (6'h26 == _T_188) begin
                                                          mem_38 <= _GEN_7;
                                                        end else begin
                                                          if (6'h26 == _T_183) begin
                                                            mem_38 <= _GEN_6;
                                                          end else begin
                                                            if (6'h26 == _T_178) begin
                                                              mem_38 <= _GEN_5;
                                                            end else begin
                                                              if (6'h26 == _T_173) begin
                                                                mem_38 <= _GEN_4;
                                                              end else begin
                                                                if (6'h26 == _T_168) begin
                                                                  mem_38 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h26 == _T_163) begin
                                                                    mem_38 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h26 == _T_158) begin
                                                                      mem_38 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h26 == _T_153) begin
                                                                        mem_38 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h27 == wPos) begin
            mem_39 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h27 == _T_308) begin
                mem_39 <= _GEN_31;
              end else begin
                if (6'h27 == _T_303) begin
                  mem_39 <= _GEN_30;
                end else begin
                  if (6'h27 == _T_298) begin
                    mem_39 <= _GEN_29;
                  end else begin
                    if (6'h27 == _T_293) begin
                      mem_39 <= _GEN_28;
                    end else begin
                      if (6'h27 == _T_288) begin
                        mem_39 <= _GEN_27;
                      end else begin
                        if (6'h27 == _T_283) begin
                          mem_39 <= _GEN_26;
                        end else begin
                          if (6'h27 == _T_278) begin
                            mem_39 <= _GEN_25;
                          end else begin
                            if (6'h27 == _T_273) begin
                              mem_39 <= _GEN_24;
                            end else begin
                              if (6'h27 == _T_268) begin
                                mem_39 <= _GEN_23;
                              end else begin
                                if (6'h27 == _T_263) begin
                                  mem_39 <= _GEN_22;
                                end else begin
                                  if (6'h27 == _T_258) begin
                                    mem_39 <= _GEN_21;
                                  end else begin
                                    if (6'h27 == _T_253) begin
                                      mem_39 <= _GEN_20;
                                    end else begin
                                      if (6'h27 == _T_248) begin
                                        mem_39 <= _GEN_19;
                                      end else begin
                                        if (6'h27 == _T_243) begin
                                          mem_39 <= _GEN_18;
                                        end else begin
                                          if (6'h27 == _T_238) begin
                                            mem_39 <= _GEN_17;
                                          end else begin
                                            if (6'h27 == _T_233) begin
                                              mem_39 <= _GEN_16;
                                            end else begin
                                              if (6'h27 == _T_228) begin
                                                mem_39 <= _GEN_15;
                                              end else begin
                                                if (6'h27 == _T_223) begin
                                                  mem_39 <= _GEN_14;
                                                end else begin
                                                  if (6'h27 == _T_218) begin
                                                    mem_39 <= _GEN_13;
                                                  end else begin
                                                    if (6'h27 == _T_213) begin
                                                      mem_39 <= _GEN_12;
                                                    end else begin
                                                      if (6'h27 == _T_208) begin
                                                        mem_39 <= _GEN_11;
                                                      end else begin
                                                        if (6'h27 == _T_203) begin
                                                          mem_39 <= _GEN_10;
                                                        end else begin
                                                          if (6'h27 == _T_198) begin
                                                            mem_39 <= _GEN_9;
                                                          end else begin
                                                            if (6'h27 == _T_193) begin
                                                              mem_39 <= _GEN_8;
                                                            end else begin
                                                              if (6'h27 == _T_188) begin
                                                                mem_39 <= _GEN_7;
                                                              end else begin
                                                                if (6'h27 == _T_183) begin
                                                                  mem_39 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h27 == _T_178) begin
                                                                    mem_39 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h27 == _T_173) begin
                                                                      mem_39 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h27 == _T_168) begin
                                                                        mem_39 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h27 == _T_163) begin
                                                                          mem_39 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h27 == _T_158) begin
                                                                            mem_39 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h27 == _T_153) begin
                                                                              mem_39 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h27 == _T_308) begin
              mem_39 <= _GEN_31;
            end else begin
              if (6'h27 == _T_303) begin
                mem_39 <= _GEN_30;
              end else begin
                if (6'h27 == _T_298) begin
                  mem_39 <= _GEN_29;
                end else begin
                  if (6'h27 == _T_293) begin
                    mem_39 <= _GEN_28;
                  end else begin
                    if (6'h27 == _T_288) begin
                      mem_39 <= _GEN_27;
                    end else begin
                      if (6'h27 == _T_283) begin
                        mem_39 <= _GEN_26;
                      end else begin
                        if (6'h27 == _T_278) begin
                          mem_39 <= _GEN_25;
                        end else begin
                          if (6'h27 == _T_273) begin
                            mem_39 <= _GEN_24;
                          end else begin
                            if (6'h27 == _T_268) begin
                              mem_39 <= _GEN_23;
                            end else begin
                              if (6'h27 == _T_263) begin
                                mem_39 <= _GEN_22;
                              end else begin
                                if (6'h27 == _T_258) begin
                                  mem_39 <= _GEN_21;
                                end else begin
                                  if (6'h27 == _T_253) begin
                                    mem_39 <= _GEN_20;
                                  end else begin
                                    if (6'h27 == _T_248) begin
                                      mem_39 <= _GEN_19;
                                    end else begin
                                      if (6'h27 == _T_243) begin
                                        mem_39 <= _GEN_18;
                                      end else begin
                                        if (6'h27 == _T_238) begin
                                          mem_39 <= _GEN_17;
                                        end else begin
                                          if (6'h27 == _T_233) begin
                                            mem_39 <= _GEN_16;
                                          end else begin
                                            if (6'h27 == _T_228) begin
                                              mem_39 <= _GEN_15;
                                            end else begin
                                              if (6'h27 == _T_223) begin
                                                mem_39 <= _GEN_14;
                                              end else begin
                                                if (6'h27 == _T_218) begin
                                                  mem_39 <= _GEN_13;
                                                end else begin
                                                  if (6'h27 == _T_213) begin
                                                    mem_39 <= _GEN_12;
                                                  end else begin
                                                    if (6'h27 == _T_208) begin
                                                      mem_39 <= _GEN_11;
                                                    end else begin
                                                      if (6'h27 == _T_203) begin
                                                        mem_39 <= _GEN_10;
                                                      end else begin
                                                        if (6'h27 == _T_198) begin
                                                          mem_39 <= _GEN_9;
                                                        end else begin
                                                          if (6'h27 == _T_193) begin
                                                            mem_39 <= _GEN_8;
                                                          end else begin
                                                            if (6'h27 == _T_188) begin
                                                              mem_39 <= _GEN_7;
                                                            end else begin
                                                              if (6'h27 == _T_183) begin
                                                                mem_39 <= _GEN_6;
                                                              end else begin
                                                                if (6'h27 == _T_178) begin
                                                                  mem_39 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h27 == _T_173) begin
                                                                    mem_39 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h27 == _T_168) begin
                                                                      mem_39 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h27 == _T_163) begin
                                                                        mem_39 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h27 == _T_158) begin
                                                                          mem_39 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h27 == _T_153) begin
                                                                            mem_39 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h27 == _T_308) begin
            mem_39 <= _GEN_31;
          end else begin
            if (6'h27 == _T_303) begin
              mem_39 <= _GEN_30;
            end else begin
              if (6'h27 == _T_298) begin
                mem_39 <= _GEN_29;
              end else begin
                if (6'h27 == _T_293) begin
                  mem_39 <= _GEN_28;
                end else begin
                  if (6'h27 == _T_288) begin
                    mem_39 <= _GEN_27;
                  end else begin
                    if (6'h27 == _T_283) begin
                      mem_39 <= _GEN_26;
                    end else begin
                      if (6'h27 == _T_278) begin
                        mem_39 <= _GEN_25;
                      end else begin
                        if (6'h27 == _T_273) begin
                          mem_39 <= _GEN_24;
                        end else begin
                          if (6'h27 == _T_268) begin
                            mem_39 <= _GEN_23;
                          end else begin
                            if (6'h27 == _T_263) begin
                              mem_39 <= _GEN_22;
                            end else begin
                              if (6'h27 == _T_258) begin
                                mem_39 <= _GEN_21;
                              end else begin
                                if (6'h27 == _T_253) begin
                                  mem_39 <= _GEN_20;
                                end else begin
                                  if (6'h27 == _T_248) begin
                                    mem_39 <= _GEN_19;
                                  end else begin
                                    if (6'h27 == _T_243) begin
                                      mem_39 <= _GEN_18;
                                    end else begin
                                      if (6'h27 == _T_238) begin
                                        mem_39 <= _GEN_17;
                                      end else begin
                                        if (6'h27 == _T_233) begin
                                          mem_39 <= _GEN_16;
                                        end else begin
                                          if (6'h27 == _T_228) begin
                                            mem_39 <= _GEN_15;
                                          end else begin
                                            if (6'h27 == _T_223) begin
                                              mem_39 <= _GEN_14;
                                            end else begin
                                              if (6'h27 == _T_218) begin
                                                mem_39 <= _GEN_13;
                                              end else begin
                                                if (6'h27 == _T_213) begin
                                                  mem_39 <= _GEN_12;
                                                end else begin
                                                  if (6'h27 == _T_208) begin
                                                    mem_39 <= _GEN_11;
                                                  end else begin
                                                    if (6'h27 == _T_203) begin
                                                      mem_39 <= _GEN_10;
                                                    end else begin
                                                      if (6'h27 == _T_198) begin
                                                        mem_39 <= _GEN_9;
                                                      end else begin
                                                        if (6'h27 == _T_193) begin
                                                          mem_39 <= _GEN_8;
                                                        end else begin
                                                          if (6'h27 == _T_188) begin
                                                            mem_39 <= _GEN_7;
                                                          end else begin
                                                            if (6'h27 == _T_183) begin
                                                              mem_39 <= _GEN_6;
                                                            end else begin
                                                              if (6'h27 == _T_178) begin
                                                                mem_39 <= _GEN_5;
                                                              end else begin
                                                                if (6'h27 == _T_173) begin
                                                                  mem_39 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h27 == _T_168) begin
                                                                    mem_39 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h27 == _T_163) begin
                                                                      mem_39 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h27 == _T_158) begin
                                                                        mem_39 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h27 == _T_153) begin
                                                                          mem_39 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h27 == _T_308) begin
          mem_39 <= _GEN_31;
        end else begin
          if (6'h27 == _T_303) begin
            mem_39 <= _GEN_30;
          end else begin
            if (6'h27 == _T_298) begin
              mem_39 <= _GEN_29;
            end else begin
              if (6'h27 == _T_293) begin
                mem_39 <= _GEN_28;
              end else begin
                if (6'h27 == _T_288) begin
                  mem_39 <= _GEN_27;
                end else begin
                  if (6'h27 == _T_283) begin
                    mem_39 <= _GEN_26;
                  end else begin
                    if (6'h27 == _T_278) begin
                      mem_39 <= _GEN_25;
                    end else begin
                      if (6'h27 == _T_273) begin
                        mem_39 <= _GEN_24;
                      end else begin
                        if (6'h27 == _T_268) begin
                          mem_39 <= _GEN_23;
                        end else begin
                          if (6'h27 == _T_263) begin
                            mem_39 <= _GEN_22;
                          end else begin
                            if (6'h27 == _T_258) begin
                              mem_39 <= _GEN_21;
                            end else begin
                              if (6'h27 == _T_253) begin
                                mem_39 <= _GEN_20;
                              end else begin
                                if (6'h27 == _T_248) begin
                                  mem_39 <= _GEN_19;
                                end else begin
                                  if (6'h27 == _T_243) begin
                                    mem_39 <= _GEN_18;
                                  end else begin
                                    if (6'h27 == _T_238) begin
                                      mem_39 <= _GEN_17;
                                    end else begin
                                      if (6'h27 == _T_233) begin
                                        mem_39 <= _GEN_16;
                                      end else begin
                                        if (6'h27 == _T_228) begin
                                          mem_39 <= _GEN_15;
                                        end else begin
                                          if (6'h27 == _T_223) begin
                                            mem_39 <= _GEN_14;
                                          end else begin
                                            if (6'h27 == _T_218) begin
                                              mem_39 <= _GEN_13;
                                            end else begin
                                              if (6'h27 == _T_213) begin
                                                mem_39 <= _GEN_12;
                                              end else begin
                                                if (6'h27 == _T_208) begin
                                                  mem_39 <= _GEN_11;
                                                end else begin
                                                  if (6'h27 == _T_203) begin
                                                    mem_39 <= _GEN_10;
                                                  end else begin
                                                    if (6'h27 == _T_198) begin
                                                      mem_39 <= _GEN_9;
                                                    end else begin
                                                      if (6'h27 == _T_193) begin
                                                        mem_39 <= _GEN_8;
                                                      end else begin
                                                        if (6'h27 == _T_188) begin
                                                          mem_39 <= _GEN_7;
                                                        end else begin
                                                          if (6'h27 == _T_183) begin
                                                            mem_39 <= _GEN_6;
                                                          end else begin
                                                            if (6'h27 == _T_178) begin
                                                              mem_39 <= _GEN_5;
                                                            end else begin
                                                              if (6'h27 == _T_173) begin
                                                                mem_39 <= _GEN_4;
                                                              end else begin
                                                                if (6'h27 == _T_168) begin
                                                                  mem_39 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h27 == _T_163) begin
                                                                    mem_39 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h27 == _T_158) begin
                                                                      mem_39 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h27 == _T_153) begin
                                                                        mem_39 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h28 == wPos) begin
            mem_40 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h28 == _T_308) begin
                mem_40 <= _GEN_31;
              end else begin
                if (6'h28 == _T_303) begin
                  mem_40 <= _GEN_30;
                end else begin
                  if (6'h28 == _T_298) begin
                    mem_40 <= _GEN_29;
                  end else begin
                    if (6'h28 == _T_293) begin
                      mem_40 <= _GEN_28;
                    end else begin
                      if (6'h28 == _T_288) begin
                        mem_40 <= _GEN_27;
                      end else begin
                        if (6'h28 == _T_283) begin
                          mem_40 <= _GEN_26;
                        end else begin
                          if (6'h28 == _T_278) begin
                            mem_40 <= _GEN_25;
                          end else begin
                            if (6'h28 == _T_273) begin
                              mem_40 <= _GEN_24;
                            end else begin
                              if (6'h28 == _T_268) begin
                                mem_40 <= _GEN_23;
                              end else begin
                                if (6'h28 == _T_263) begin
                                  mem_40 <= _GEN_22;
                                end else begin
                                  if (6'h28 == _T_258) begin
                                    mem_40 <= _GEN_21;
                                  end else begin
                                    if (6'h28 == _T_253) begin
                                      mem_40 <= _GEN_20;
                                    end else begin
                                      if (6'h28 == _T_248) begin
                                        mem_40 <= _GEN_19;
                                      end else begin
                                        if (6'h28 == _T_243) begin
                                          mem_40 <= _GEN_18;
                                        end else begin
                                          if (6'h28 == _T_238) begin
                                            mem_40 <= _GEN_17;
                                          end else begin
                                            if (6'h28 == _T_233) begin
                                              mem_40 <= _GEN_16;
                                            end else begin
                                              if (6'h28 == _T_228) begin
                                                mem_40 <= _GEN_15;
                                              end else begin
                                                if (6'h28 == _T_223) begin
                                                  mem_40 <= _GEN_14;
                                                end else begin
                                                  if (6'h28 == _T_218) begin
                                                    mem_40 <= _GEN_13;
                                                  end else begin
                                                    if (6'h28 == _T_213) begin
                                                      mem_40 <= _GEN_12;
                                                    end else begin
                                                      if (6'h28 == _T_208) begin
                                                        mem_40 <= _GEN_11;
                                                      end else begin
                                                        if (6'h28 == _T_203) begin
                                                          mem_40 <= _GEN_10;
                                                        end else begin
                                                          if (6'h28 == _T_198) begin
                                                            mem_40 <= _GEN_9;
                                                          end else begin
                                                            if (6'h28 == _T_193) begin
                                                              mem_40 <= _GEN_8;
                                                            end else begin
                                                              if (6'h28 == _T_188) begin
                                                                mem_40 <= _GEN_7;
                                                              end else begin
                                                                if (6'h28 == _T_183) begin
                                                                  mem_40 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h28 == _T_178) begin
                                                                    mem_40 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h28 == _T_173) begin
                                                                      mem_40 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h28 == _T_168) begin
                                                                        mem_40 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h28 == _T_163) begin
                                                                          mem_40 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h28 == _T_158) begin
                                                                            mem_40 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h28 == _T_153) begin
                                                                              mem_40 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h28 == _T_308) begin
              mem_40 <= _GEN_31;
            end else begin
              if (6'h28 == _T_303) begin
                mem_40 <= _GEN_30;
              end else begin
                if (6'h28 == _T_298) begin
                  mem_40 <= _GEN_29;
                end else begin
                  if (6'h28 == _T_293) begin
                    mem_40 <= _GEN_28;
                  end else begin
                    if (6'h28 == _T_288) begin
                      mem_40 <= _GEN_27;
                    end else begin
                      if (6'h28 == _T_283) begin
                        mem_40 <= _GEN_26;
                      end else begin
                        if (6'h28 == _T_278) begin
                          mem_40 <= _GEN_25;
                        end else begin
                          if (6'h28 == _T_273) begin
                            mem_40 <= _GEN_24;
                          end else begin
                            if (6'h28 == _T_268) begin
                              mem_40 <= _GEN_23;
                            end else begin
                              if (6'h28 == _T_263) begin
                                mem_40 <= _GEN_22;
                              end else begin
                                if (6'h28 == _T_258) begin
                                  mem_40 <= _GEN_21;
                                end else begin
                                  if (6'h28 == _T_253) begin
                                    mem_40 <= _GEN_20;
                                  end else begin
                                    if (6'h28 == _T_248) begin
                                      mem_40 <= _GEN_19;
                                    end else begin
                                      if (6'h28 == _T_243) begin
                                        mem_40 <= _GEN_18;
                                      end else begin
                                        if (6'h28 == _T_238) begin
                                          mem_40 <= _GEN_17;
                                        end else begin
                                          if (6'h28 == _T_233) begin
                                            mem_40 <= _GEN_16;
                                          end else begin
                                            if (6'h28 == _T_228) begin
                                              mem_40 <= _GEN_15;
                                            end else begin
                                              if (6'h28 == _T_223) begin
                                                mem_40 <= _GEN_14;
                                              end else begin
                                                if (6'h28 == _T_218) begin
                                                  mem_40 <= _GEN_13;
                                                end else begin
                                                  if (6'h28 == _T_213) begin
                                                    mem_40 <= _GEN_12;
                                                  end else begin
                                                    if (6'h28 == _T_208) begin
                                                      mem_40 <= _GEN_11;
                                                    end else begin
                                                      if (6'h28 == _T_203) begin
                                                        mem_40 <= _GEN_10;
                                                      end else begin
                                                        if (6'h28 == _T_198) begin
                                                          mem_40 <= _GEN_9;
                                                        end else begin
                                                          if (6'h28 == _T_193) begin
                                                            mem_40 <= _GEN_8;
                                                          end else begin
                                                            if (6'h28 == _T_188) begin
                                                              mem_40 <= _GEN_7;
                                                            end else begin
                                                              if (6'h28 == _T_183) begin
                                                                mem_40 <= _GEN_6;
                                                              end else begin
                                                                if (6'h28 == _T_178) begin
                                                                  mem_40 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h28 == _T_173) begin
                                                                    mem_40 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h28 == _T_168) begin
                                                                      mem_40 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h28 == _T_163) begin
                                                                        mem_40 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h28 == _T_158) begin
                                                                          mem_40 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h28 == _T_153) begin
                                                                            mem_40 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h28 == _T_308) begin
            mem_40 <= _GEN_31;
          end else begin
            if (6'h28 == _T_303) begin
              mem_40 <= _GEN_30;
            end else begin
              if (6'h28 == _T_298) begin
                mem_40 <= _GEN_29;
              end else begin
                if (6'h28 == _T_293) begin
                  mem_40 <= _GEN_28;
                end else begin
                  if (6'h28 == _T_288) begin
                    mem_40 <= _GEN_27;
                  end else begin
                    if (6'h28 == _T_283) begin
                      mem_40 <= _GEN_26;
                    end else begin
                      if (6'h28 == _T_278) begin
                        mem_40 <= _GEN_25;
                      end else begin
                        if (6'h28 == _T_273) begin
                          mem_40 <= _GEN_24;
                        end else begin
                          if (6'h28 == _T_268) begin
                            mem_40 <= _GEN_23;
                          end else begin
                            if (6'h28 == _T_263) begin
                              mem_40 <= _GEN_22;
                            end else begin
                              if (6'h28 == _T_258) begin
                                mem_40 <= _GEN_21;
                              end else begin
                                if (6'h28 == _T_253) begin
                                  mem_40 <= _GEN_20;
                                end else begin
                                  if (6'h28 == _T_248) begin
                                    mem_40 <= _GEN_19;
                                  end else begin
                                    if (6'h28 == _T_243) begin
                                      mem_40 <= _GEN_18;
                                    end else begin
                                      if (6'h28 == _T_238) begin
                                        mem_40 <= _GEN_17;
                                      end else begin
                                        if (6'h28 == _T_233) begin
                                          mem_40 <= _GEN_16;
                                        end else begin
                                          if (6'h28 == _T_228) begin
                                            mem_40 <= _GEN_15;
                                          end else begin
                                            if (6'h28 == _T_223) begin
                                              mem_40 <= _GEN_14;
                                            end else begin
                                              if (6'h28 == _T_218) begin
                                                mem_40 <= _GEN_13;
                                              end else begin
                                                if (6'h28 == _T_213) begin
                                                  mem_40 <= _GEN_12;
                                                end else begin
                                                  if (6'h28 == _T_208) begin
                                                    mem_40 <= _GEN_11;
                                                  end else begin
                                                    if (6'h28 == _T_203) begin
                                                      mem_40 <= _GEN_10;
                                                    end else begin
                                                      if (6'h28 == _T_198) begin
                                                        mem_40 <= _GEN_9;
                                                      end else begin
                                                        if (6'h28 == _T_193) begin
                                                          mem_40 <= _GEN_8;
                                                        end else begin
                                                          if (6'h28 == _T_188) begin
                                                            mem_40 <= _GEN_7;
                                                          end else begin
                                                            if (6'h28 == _T_183) begin
                                                              mem_40 <= _GEN_6;
                                                            end else begin
                                                              if (6'h28 == _T_178) begin
                                                                mem_40 <= _GEN_5;
                                                              end else begin
                                                                if (6'h28 == _T_173) begin
                                                                  mem_40 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h28 == _T_168) begin
                                                                    mem_40 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h28 == _T_163) begin
                                                                      mem_40 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h28 == _T_158) begin
                                                                        mem_40 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h28 == _T_153) begin
                                                                          mem_40 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h28 == _T_308) begin
          mem_40 <= _GEN_31;
        end else begin
          if (6'h28 == _T_303) begin
            mem_40 <= _GEN_30;
          end else begin
            if (6'h28 == _T_298) begin
              mem_40 <= _GEN_29;
            end else begin
              if (6'h28 == _T_293) begin
                mem_40 <= _GEN_28;
              end else begin
                if (6'h28 == _T_288) begin
                  mem_40 <= _GEN_27;
                end else begin
                  if (6'h28 == _T_283) begin
                    mem_40 <= _GEN_26;
                  end else begin
                    if (6'h28 == _T_278) begin
                      mem_40 <= _GEN_25;
                    end else begin
                      if (6'h28 == _T_273) begin
                        mem_40 <= _GEN_24;
                      end else begin
                        if (6'h28 == _T_268) begin
                          mem_40 <= _GEN_23;
                        end else begin
                          if (6'h28 == _T_263) begin
                            mem_40 <= _GEN_22;
                          end else begin
                            if (6'h28 == _T_258) begin
                              mem_40 <= _GEN_21;
                            end else begin
                              if (6'h28 == _T_253) begin
                                mem_40 <= _GEN_20;
                              end else begin
                                if (6'h28 == _T_248) begin
                                  mem_40 <= _GEN_19;
                                end else begin
                                  if (6'h28 == _T_243) begin
                                    mem_40 <= _GEN_18;
                                  end else begin
                                    if (6'h28 == _T_238) begin
                                      mem_40 <= _GEN_17;
                                    end else begin
                                      if (6'h28 == _T_233) begin
                                        mem_40 <= _GEN_16;
                                      end else begin
                                        if (6'h28 == _T_228) begin
                                          mem_40 <= _GEN_15;
                                        end else begin
                                          if (6'h28 == _T_223) begin
                                            mem_40 <= _GEN_14;
                                          end else begin
                                            if (6'h28 == _T_218) begin
                                              mem_40 <= _GEN_13;
                                            end else begin
                                              if (6'h28 == _T_213) begin
                                                mem_40 <= _GEN_12;
                                              end else begin
                                                if (6'h28 == _T_208) begin
                                                  mem_40 <= _GEN_11;
                                                end else begin
                                                  if (6'h28 == _T_203) begin
                                                    mem_40 <= _GEN_10;
                                                  end else begin
                                                    if (6'h28 == _T_198) begin
                                                      mem_40 <= _GEN_9;
                                                    end else begin
                                                      if (6'h28 == _T_193) begin
                                                        mem_40 <= _GEN_8;
                                                      end else begin
                                                        if (6'h28 == _T_188) begin
                                                          mem_40 <= _GEN_7;
                                                        end else begin
                                                          if (6'h28 == _T_183) begin
                                                            mem_40 <= _GEN_6;
                                                          end else begin
                                                            if (6'h28 == _T_178) begin
                                                              mem_40 <= _GEN_5;
                                                            end else begin
                                                              if (6'h28 == _T_173) begin
                                                                mem_40 <= _GEN_4;
                                                              end else begin
                                                                if (6'h28 == _T_168) begin
                                                                  mem_40 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h28 == _T_163) begin
                                                                    mem_40 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h28 == _T_158) begin
                                                                      mem_40 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h28 == _T_153) begin
                                                                        mem_40 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h29 == wPos) begin
            mem_41 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h29 == _T_308) begin
                mem_41 <= _GEN_31;
              end else begin
                if (6'h29 == _T_303) begin
                  mem_41 <= _GEN_30;
                end else begin
                  if (6'h29 == _T_298) begin
                    mem_41 <= _GEN_29;
                  end else begin
                    if (6'h29 == _T_293) begin
                      mem_41 <= _GEN_28;
                    end else begin
                      if (6'h29 == _T_288) begin
                        mem_41 <= _GEN_27;
                      end else begin
                        if (6'h29 == _T_283) begin
                          mem_41 <= _GEN_26;
                        end else begin
                          if (6'h29 == _T_278) begin
                            mem_41 <= _GEN_25;
                          end else begin
                            if (6'h29 == _T_273) begin
                              mem_41 <= _GEN_24;
                            end else begin
                              if (6'h29 == _T_268) begin
                                mem_41 <= _GEN_23;
                              end else begin
                                if (6'h29 == _T_263) begin
                                  mem_41 <= _GEN_22;
                                end else begin
                                  if (6'h29 == _T_258) begin
                                    mem_41 <= _GEN_21;
                                  end else begin
                                    if (6'h29 == _T_253) begin
                                      mem_41 <= _GEN_20;
                                    end else begin
                                      if (6'h29 == _T_248) begin
                                        mem_41 <= _GEN_19;
                                      end else begin
                                        if (6'h29 == _T_243) begin
                                          mem_41 <= _GEN_18;
                                        end else begin
                                          if (6'h29 == _T_238) begin
                                            mem_41 <= _GEN_17;
                                          end else begin
                                            if (6'h29 == _T_233) begin
                                              mem_41 <= _GEN_16;
                                            end else begin
                                              if (6'h29 == _T_228) begin
                                                mem_41 <= _GEN_15;
                                              end else begin
                                                if (6'h29 == _T_223) begin
                                                  mem_41 <= _GEN_14;
                                                end else begin
                                                  if (6'h29 == _T_218) begin
                                                    mem_41 <= _GEN_13;
                                                  end else begin
                                                    if (6'h29 == _T_213) begin
                                                      mem_41 <= _GEN_12;
                                                    end else begin
                                                      if (6'h29 == _T_208) begin
                                                        mem_41 <= _GEN_11;
                                                      end else begin
                                                        if (6'h29 == _T_203) begin
                                                          mem_41 <= _GEN_10;
                                                        end else begin
                                                          if (6'h29 == _T_198) begin
                                                            mem_41 <= _GEN_9;
                                                          end else begin
                                                            if (6'h29 == _T_193) begin
                                                              mem_41 <= _GEN_8;
                                                            end else begin
                                                              if (6'h29 == _T_188) begin
                                                                mem_41 <= _GEN_7;
                                                              end else begin
                                                                if (6'h29 == _T_183) begin
                                                                  mem_41 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h29 == _T_178) begin
                                                                    mem_41 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h29 == _T_173) begin
                                                                      mem_41 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h29 == _T_168) begin
                                                                        mem_41 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h29 == _T_163) begin
                                                                          mem_41 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h29 == _T_158) begin
                                                                            mem_41 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h29 == _T_153) begin
                                                                              mem_41 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h29 == _T_308) begin
              mem_41 <= _GEN_31;
            end else begin
              if (6'h29 == _T_303) begin
                mem_41 <= _GEN_30;
              end else begin
                if (6'h29 == _T_298) begin
                  mem_41 <= _GEN_29;
                end else begin
                  if (6'h29 == _T_293) begin
                    mem_41 <= _GEN_28;
                  end else begin
                    if (6'h29 == _T_288) begin
                      mem_41 <= _GEN_27;
                    end else begin
                      if (6'h29 == _T_283) begin
                        mem_41 <= _GEN_26;
                      end else begin
                        if (6'h29 == _T_278) begin
                          mem_41 <= _GEN_25;
                        end else begin
                          if (6'h29 == _T_273) begin
                            mem_41 <= _GEN_24;
                          end else begin
                            if (6'h29 == _T_268) begin
                              mem_41 <= _GEN_23;
                            end else begin
                              if (6'h29 == _T_263) begin
                                mem_41 <= _GEN_22;
                              end else begin
                                if (6'h29 == _T_258) begin
                                  mem_41 <= _GEN_21;
                                end else begin
                                  if (6'h29 == _T_253) begin
                                    mem_41 <= _GEN_20;
                                  end else begin
                                    if (6'h29 == _T_248) begin
                                      mem_41 <= _GEN_19;
                                    end else begin
                                      if (6'h29 == _T_243) begin
                                        mem_41 <= _GEN_18;
                                      end else begin
                                        if (6'h29 == _T_238) begin
                                          mem_41 <= _GEN_17;
                                        end else begin
                                          if (6'h29 == _T_233) begin
                                            mem_41 <= _GEN_16;
                                          end else begin
                                            if (6'h29 == _T_228) begin
                                              mem_41 <= _GEN_15;
                                            end else begin
                                              if (6'h29 == _T_223) begin
                                                mem_41 <= _GEN_14;
                                              end else begin
                                                if (6'h29 == _T_218) begin
                                                  mem_41 <= _GEN_13;
                                                end else begin
                                                  if (6'h29 == _T_213) begin
                                                    mem_41 <= _GEN_12;
                                                  end else begin
                                                    if (6'h29 == _T_208) begin
                                                      mem_41 <= _GEN_11;
                                                    end else begin
                                                      if (6'h29 == _T_203) begin
                                                        mem_41 <= _GEN_10;
                                                      end else begin
                                                        if (6'h29 == _T_198) begin
                                                          mem_41 <= _GEN_9;
                                                        end else begin
                                                          if (6'h29 == _T_193) begin
                                                            mem_41 <= _GEN_8;
                                                          end else begin
                                                            if (6'h29 == _T_188) begin
                                                              mem_41 <= _GEN_7;
                                                            end else begin
                                                              if (6'h29 == _T_183) begin
                                                                mem_41 <= _GEN_6;
                                                              end else begin
                                                                if (6'h29 == _T_178) begin
                                                                  mem_41 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h29 == _T_173) begin
                                                                    mem_41 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h29 == _T_168) begin
                                                                      mem_41 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h29 == _T_163) begin
                                                                        mem_41 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h29 == _T_158) begin
                                                                          mem_41 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h29 == _T_153) begin
                                                                            mem_41 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h29 == _T_308) begin
            mem_41 <= _GEN_31;
          end else begin
            if (6'h29 == _T_303) begin
              mem_41 <= _GEN_30;
            end else begin
              if (6'h29 == _T_298) begin
                mem_41 <= _GEN_29;
              end else begin
                if (6'h29 == _T_293) begin
                  mem_41 <= _GEN_28;
                end else begin
                  if (6'h29 == _T_288) begin
                    mem_41 <= _GEN_27;
                  end else begin
                    if (6'h29 == _T_283) begin
                      mem_41 <= _GEN_26;
                    end else begin
                      if (6'h29 == _T_278) begin
                        mem_41 <= _GEN_25;
                      end else begin
                        if (6'h29 == _T_273) begin
                          mem_41 <= _GEN_24;
                        end else begin
                          if (6'h29 == _T_268) begin
                            mem_41 <= _GEN_23;
                          end else begin
                            if (6'h29 == _T_263) begin
                              mem_41 <= _GEN_22;
                            end else begin
                              if (6'h29 == _T_258) begin
                                mem_41 <= _GEN_21;
                              end else begin
                                if (6'h29 == _T_253) begin
                                  mem_41 <= _GEN_20;
                                end else begin
                                  if (6'h29 == _T_248) begin
                                    mem_41 <= _GEN_19;
                                  end else begin
                                    if (6'h29 == _T_243) begin
                                      mem_41 <= _GEN_18;
                                    end else begin
                                      if (6'h29 == _T_238) begin
                                        mem_41 <= _GEN_17;
                                      end else begin
                                        if (6'h29 == _T_233) begin
                                          mem_41 <= _GEN_16;
                                        end else begin
                                          if (6'h29 == _T_228) begin
                                            mem_41 <= _GEN_15;
                                          end else begin
                                            if (6'h29 == _T_223) begin
                                              mem_41 <= _GEN_14;
                                            end else begin
                                              if (6'h29 == _T_218) begin
                                                mem_41 <= _GEN_13;
                                              end else begin
                                                if (6'h29 == _T_213) begin
                                                  mem_41 <= _GEN_12;
                                                end else begin
                                                  if (6'h29 == _T_208) begin
                                                    mem_41 <= _GEN_11;
                                                  end else begin
                                                    if (6'h29 == _T_203) begin
                                                      mem_41 <= _GEN_10;
                                                    end else begin
                                                      if (6'h29 == _T_198) begin
                                                        mem_41 <= _GEN_9;
                                                      end else begin
                                                        if (6'h29 == _T_193) begin
                                                          mem_41 <= _GEN_8;
                                                        end else begin
                                                          if (6'h29 == _T_188) begin
                                                            mem_41 <= _GEN_7;
                                                          end else begin
                                                            if (6'h29 == _T_183) begin
                                                              mem_41 <= _GEN_6;
                                                            end else begin
                                                              if (6'h29 == _T_178) begin
                                                                mem_41 <= _GEN_5;
                                                              end else begin
                                                                if (6'h29 == _T_173) begin
                                                                  mem_41 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h29 == _T_168) begin
                                                                    mem_41 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h29 == _T_163) begin
                                                                      mem_41 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h29 == _T_158) begin
                                                                        mem_41 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h29 == _T_153) begin
                                                                          mem_41 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h29 == _T_308) begin
          mem_41 <= _GEN_31;
        end else begin
          if (6'h29 == _T_303) begin
            mem_41 <= _GEN_30;
          end else begin
            if (6'h29 == _T_298) begin
              mem_41 <= _GEN_29;
            end else begin
              if (6'h29 == _T_293) begin
                mem_41 <= _GEN_28;
              end else begin
                if (6'h29 == _T_288) begin
                  mem_41 <= _GEN_27;
                end else begin
                  if (6'h29 == _T_283) begin
                    mem_41 <= _GEN_26;
                  end else begin
                    if (6'h29 == _T_278) begin
                      mem_41 <= _GEN_25;
                    end else begin
                      if (6'h29 == _T_273) begin
                        mem_41 <= _GEN_24;
                      end else begin
                        if (6'h29 == _T_268) begin
                          mem_41 <= _GEN_23;
                        end else begin
                          if (6'h29 == _T_263) begin
                            mem_41 <= _GEN_22;
                          end else begin
                            if (6'h29 == _T_258) begin
                              mem_41 <= _GEN_21;
                            end else begin
                              if (6'h29 == _T_253) begin
                                mem_41 <= _GEN_20;
                              end else begin
                                if (6'h29 == _T_248) begin
                                  mem_41 <= _GEN_19;
                                end else begin
                                  if (6'h29 == _T_243) begin
                                    mem_41 <= _GEN_18;
                                  end else begin
                                    if (6'h29 == _T_238) begin
                                      mem_41 <= _GEN_17;
                                    end else begin
                                      if (6'h29 == _T_233) begin
                                        mem_41 <= _GEN_16;
                                      end else begin
                                        if (6'h29 == _T_228) begin
                                          mem_41 <= _GEN_15;
                                        end else begin
                                          if (6'h29 == _T_223) begin
                                            mem_41 <= _GEN_14;
                                          end else begin
                                            if (6'h29 == _T_218) begin
                                              mem_41 <= _GEN_13;
                                            end else begin
                                              if (6'h29 == _T_213) begin
                                                mem_41 <= _GEN_12;
                                              end else begin
                                                if (6'h29 == _T_208) begin
                                                  mem_41 <= _GEN_11;
                                                end else begin
                                                  if (6'h29 == _T_203) begin
                                                    mem_41 <= _GEN_10;
                                                  end else begin
                                                    if (6'h29 == _T_198) begin
                                                      mem_41 <= _GEN_9;
                                                    end else begin
                                                      if (6'h29 == _T_193) begin
                                                        mem_41 <= _GEN_8;
                                                      end else begin
                                                        if (6'h29 == _T_188) begin
                                                          mem_41 <= _GEN_7;
                                                        end else begin
                                                          if (6'h29 == _T_183) begin
                                                            mem_41 <= _GEN_6;
                                                          end else begin
                                                            if (6'h29 == _T_178) begin
                                                              mem_41 <= _GEN_5;
                                                            end else begin
                                                              if (6'h29 == _T_173) begin
                                                                mem_41 <= _GEN_4;
                                                              end else begin
                                                                if (6'h29 == _T_168) begin
                                                                  mem_41 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h29 == _T_163) begin
                                                                    mem_41 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h29 == _T_158) begin
                                                                      mem_41 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h29 == _T_153) begin
                                                                        mem_41 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h2a == wPos) begin
            mem_42 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h2a == _T_308) begin
                mem_42 <= _GEN_31;
              end else begin
                if (6'h2a == _T_303) begin
                  mem_42 <= _GEN_30;
                end else begin
                  if (6'h2a == _T_298) begin
                    mem_42 <= _GEN_29;
                  end else begin
                    if (6'h2a == _T_293) begin
                      mem_42 <= _GEN_28;
                    end else begin
                      if (6'h2a == _T_288) begin
                        mem_42 <= _GEN_27;
                      end else begin
                        if (6'h2a == _T_283) begin
                          mem_42 <= _GEN_26;
                        end else begin
                          if (6'h2a == _T_278) begin
                            mem_42 <= _GEN_25;
                          end else begin
                            if (6'h2a == _T_273) begin
                              mem_42 <= _GEN_24;
                            end else begin
                              if (6'h2a == _T_268) begin
                                mem_42 <= _GEN_23;
                              end else begin
                                if (6'h2a == _T_263) begin
                                  mem_42 <= _GEN_22;
                                end else begin
                                  if (6'h2a == _T_258) begin
                                    mem_42 <= _GEN_21;
                                  end else begin
                                    if (6'h2a == _T_253) begin
                                      mem_42 <= _GEN_20;
                                    end else begin
                                      if (6'h2a == _T_248) begin
                                        mem_42 <= _GEN_19;
                                      end else begin
                                        if (6'h2a == _T_243) begin
                                          mem_42 <= _GEN_18;
                                        end else begin
                                          if (6'h2a == _T_238) begin
                                            mem_42 <= _GEN_17;
                                          end else begin
                                            if (6'h2a == _T_233) begin
                                              mem_42 <= _GEN_16;
                                            end else begin
                                              if (6'h2a == _T_228) begin
                                                mem_42 <= _GEN_15;
                                              end else begin
                                                if (6'h2a == _T_223) begin
                                                  mem_42 <= _GEN_14;
                                                end else begin
                                                  if (6'h2a == _T_218) begin
                                                    mem_42 <= _GEN_13;
                                                  end else begin
                                                    if (6'h2a == _T_213) begin
                                                      mem_42 <= _GEN_12;
                                                    end else begin
                                                      if (6'h2a == _T_208) begin
                                                        mem_42 <= _GEN_11;
                                                      end else begin
                                                        if (6'h2a == _T_203) begin
                                                          mem_42 <= _GEN_10;
                                                        end else begin
                                                          if (6'h2a == _T_198) begin
                                                            mem_42 <= _GEN_9;
                                                          end else begin
                                                            if (6'h2a == _T_193) begin
                                                              mem_42 <= _GEN_8;
                                                            end else begin
                                                              if (6'h2a == _T_188) begin
                                                                mem_42 <= _GEN_7;
                                                              end else begin
                                                                if (6'h2a == _T_183) begin
                                                                  mem_42 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h2a == _T_178) begin
                                                                    mem_42 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h2a == _T_173) begin
                                                                      mem_42 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h2a == _T_168) begin
                                                                        mem_42 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h2a == _T_163) begin
                                                                          mem_42 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h2a == _T_158) begin
                                                                            mem_42 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h2a == _T_153) begin
                                                                              mem_42 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h2a == _T_308) begin
              mem_42 <= _GEN_31;
            end else begin
              if (6'h2a == _T_303) begin
                mem_42 <= _GEN_30;
              end else begin
                if (6'h2a == _T_298) begin
                  mem_42 <= _GEN_29;
                end else begin
                  if (6'h2a == _T_293) begin
                    mem_42 <= _GEN_28;
                  end else begin
                    if (6'h2a == _T_288) begin
                      mem_42 <= _GEN_27;
                    end else begin
                      if (6'h2a == _T_283) begin
                        mem_42 <= _GEN_26;
                      end else begin
                        if (6'h2a == _T_278) begin
                          mem_42 <= _GEN_25;
                        end else begin
                          if (6'h2a == _T_273) begin
                            mem_42 <= _GEN_24;
                          end else begin
                            if (6'h2a == _T_268) begin
                              mem_42 <= _GEN_23;
                            end else begin
                              if (6'h2a == _T_263) begin
                                mem_42 <= _GEN_22;
                              end else begin
                                if (6'h2a == _T_258) begin
                                  mem_42 <= _GEN_21;
                                end else begin
                                  if (6'h2a == _T_253) begin
                                    mem_42 <= _GEN_20;
                                  end else begin
                                    if (6'h2a == _T_248) begin
                                      mem_42 <= _GEN_19;
                                    end else begin
                                      if (6'h2a == _T_243) begin
                                        mem_42 <= _GEN_18;
                                      end else begin
                                        if (6'h2a == _T_238) begin
                                          mem_42 <= _GEN_17;
                                        end else begin
                                          if (6'h2a == _T_233) begin
                                            mem_42 <= _GEN_16;
                                          end else begin
                                            if (6'h2a == _T_228) begin
                                              mem_42 <= _GEN_15;
                                            end else begin
                                              if (6'h2a == _T_223) begin
                                                mem_42 <= _GEN_14;
                                              end else begin
                                                if (6'h2a == _T_218) begin
                                                  mem_42 <= _GEN_13;
                                                end else begin
                                                  if (6'h2a == _T_213) begin
                                                    mem_42 <= _GEN_12;
                                                  end else begin
                                                    if (6'h2a == _T_208) begin
                                                      mem_42 <= _GEN_11;
                                                    end else begin
                                                      if (6'h2a == _T_203) begin
                                                        mem_42 <= _GEN_10;
                                                      end else begin
                                                        if (6'h2a == _T_198) begin
                                                          mem_42 <= _GEN_9;
                                                        end else begin
                                                          if (6'h2a == _T_193) begin
                                                            mem_42 <= _GEN_8;
                                                          end else begin
                                                            if (6'h2a == _T_188) begin
                                                              mem_42 <= _GEN_7;
                                                            end else begin
                                                              if (6'h2a == _T_183) begin
                                                                mem_42 <= _GEN_6;
                                                              end else begin
                                                                if (6'h2a == _T_178) begin
                                                                  mem_42 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h2a == _T_173) begin
                                                                    mem_42 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h2a == _T_168) begin
                                                                      mem_42 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h2a == _T_163) begin
                                                                        mem_42 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h2a == _T_158) begin
                                                                          mem_42 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h2a == _T_153) begin
                                                                            mem_42 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h2a == _T_308) begin
            mem_42 <= _GEN_31;
          end else begin
            if (6'h2a == _T_303) begin
              mem_42 <= _GEN_30;
            end else begin
              if (6'h2a == _T_298) begin
                mem_42 <= _GEN_29;
              end else begin
                if (6'h2a == _T_293) begin
                  mem_42 <= _GEN_28;
                end else begin
                  if (6'h2a == _T_288) begin
                    mem_42 <= _GEN_27;
                  end else begin
                    if (6'h2a == _T_283) begin
                      mem_42 <= _GEN_26;
                    end else begin
                      if (6'h2a == _T_278) begin
                        mem_42 <= _GEN_25;
                      end else begin
                        if (6'h2a == _T_273) begin
                          mem_42 <= _GEN_24;
                        end else begin
                          if (6'h2a == _T_268) begin
                            mem_42 <= _GEN_23;
                          end else begin
                            if (6'h2a == _T_263) begin
                              mem_42 <= _GEN_22;
                            end else begin
                              if (6'h2a == _T_258) begin
                                mem_42 <= _GEN_21;
                              end else begin
                                if (6'h2a == _T_253) begin
                                  mem_42 <= _GEN_20;
                                end else begin
                                  if (6'h2a == _T_248) begin
                                    mem_42 <= _GEN_19;
                                  end else begin
                                    if (6'h2a == _T_243) begin
                                      mem_42 <= _GEN_18;
                                    end else begin
                                      if (6'h2a == _T_238) begin
                                        mem_42 <= _GEN_17;
                                      end else begin
                                        if (6'h2a == _T_233) begin
                                          mem_42 <= _GEN_16;
                                        end else begin
                                          if (6'h2a == _T_228) begin
                                            mem_42 <= _GEN_15;
                                          end else begin
                                            if (6'h2a == _T_223) begin
                                              mem_42 <= _GEN_14;
                                            end else begin
                                              if (6'h2a == _T_218) begin
                                                mem_42 <= _GEN_13;
                                              end else begin
                                                if (6'h2a == _T_213) begin
                                                  mem_42 <= _GEN_12;
                                                end else begin
                                                  if (6'h2a == _T_208) begin
                                                    mem_42 <= _GEN_11;
                                                  end else begin
                                                    if (6'h2a == _T_203) begin
                                                      mem_42 <= _GEN_10;
                                                    end else begin
                                                      if (6'h2a == _T_198) begin
                                                        mem_42 <= _GEN_9;
                                                      end else begin
                                                        if (6'h2a == _T_193) begin
                                                          mem_42 <= _GEN_8;
                                                        end else begin
                                                          if (6'h2a == _T_188) begin
                                                            mem_42 <= _GEN_7;
                                                          end else begin
                                                            if (6'h2a == _T_183) begin
                                                              mem_42 <= _GEN_6;
                                                            end else begin
                                                              if (6'h2a == _T_178) begin
                                                                mem_42 <= _GEN_5;
                                                              end else begin
                                                                if (6'h2a == _T_173) begin
                                                                  mem_42 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h2a == _T_168) begin
                                                                    mem_42 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h2a == _T_163) begin
                                                                      mem_42 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h2a == _T_158) begin
                                                                        mem_42 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h2a == _T_153) begin
                                                                          mem_42 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h2a == _T_308) begin
          mem_42 <= _GEN_31;
        end else begin
          if (6'h2a == _T_303) begin
            mem_42 <= _GEN_30;
          end else begin
            if (6'h2a == _T_298) begin
              mem_42 <= _GEN_29;
            end else begin
              if (6'h2a == _T_293) begin
                mem_42 <= _GEN_28;
              end else begin
                if (6'h2a == _T_288) begin
                  mem_42 <= _GEN_27;
                end else begin
                  if (6'h2a == _T_283) begin
                    mem_42 <= _GEN_26;
                  end else begin
                    if (6'h2a == _T_278) begin
                      mem_42 <= _GEN_25;
                    end else begin
                      if (6'h2a == _T_273) begin
                        mem_42 <= _GEN_24;
                      end else begin
                        if (6'h2a == _T_268) begin
                          mem_42 <= _GEN_23;
                        end else begin
                          if (6'h2a == _T_263) begin
                            mem_42 <= _GEN_22;
                          end else begin
                            if (6'h2a == _T_258) begin
                              mem_42 <= _GEN_21;
                            end else begin
                              if (6'h2a == _T_253) begin
                                mem_42 <= _GEN_20;
                              end else begin
                                if (6'h2a == _T_248) begin
                                  mem_42 <= _GEN_19;
                                end else begin
                                  if (6'h2a == _T_243) begin
                                    mem_42 <= _GEN_18;
                                  end else begin
                                    if (6'h2a == _T_238) begin
                                      mem_42 <= _GEN_17;
                                    end else begin
                                      if (6'h2a == _T_233) begin
                                        mem_42 <= _GEN_16;
                                      end else begin
                                        if (6'h2a == _T_228) begin
                                          mem_42 <= _GEN_15;
                                        end else begin
                                          if (6'h2a == _T_223) begin
                                            mem_42 <= _GEN_14;
                                          end else begin
                                            if (6'h2a == _T_218) begin
                                              mem_42 <= _GEN_13;
                                            end else begin
                                              if (6'h2a == _T_213) begin
                                                mem_42 <= _GEN_12;
                                              end else begin
                                                if (6'h2a == _T_208) begin
                                                  mem_42 <= _GEN_11;
                                                end else begin
                                                  if (6'h2a == _T_203) begin
                                                    mem_42 <= _GEN_10;
                                                  end else begin
                                                    if (6'h2a == _T_198) begin
                                                      mem_42 <= _GEN_9;
                                                    end else begin
                                                      if (6'h2a == _T_193) begin
                                                        mem_42 <= _GEN_8;
                                                      end else begin
                                                        if (6'h2a == _T_188) begin
                                                          mem_42 <= _GEN_7;
                                                        end else begin
                                                          if (6'h2a == _T_183) begin
                                                            mem_42 <= _GEN_6;
                                                          end else begin
                                                            if (6'h2a == _T_178) begin
                                                              mem_42 <= _GEN_5;
                                                            end else begin
                                                              if (6'h2a == _T_173) begin
                                                                mem_42 <= _GEN_4;
                                                              end else begin
                                                                if (6'h2a == _T_168) begin
                                                                  mem_42 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h2a == _T_163) begin
                                                                    mem_42 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h2a == _T_158) begin
                                                                      mem_42 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h2a == _T_153) begin
                                                                        mem_42 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h2b == wPos) begin
            mem_43 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h2b == _T_308) begin
                mem_43 <= _GEN_31;
              end else begin
                if (6'h2b == _T_303) begin
                  mem_43 <= _GEN_30;
                end else begin
                  if (6'h2b == _T_298) begin
                    mem_43 <= _GEN_29;
                  end else begin
                    if (6'h2b == _T_293) begin
                      mem_43 <= _GEN_28;
                    end else begin
                      if (6'h2b == _T_288) begin
                        mem_43 <= _GEN_27;
                      end else begin
                        if (6'h2b == _T_283) begin
                          mem_43 <= _GEN_26;
                        end else begin
                          if (6'h2b == _T_278) begin
                            mem_43 <= _GEN_25;
                          end else begin
                            if (6'h2b == _T_273) begin
                              mem_43 <= _GEN_24;
                            end else begin
                              if (6'h2b == _T_268) begin
                                mem_43 <= _GEN_23;
                              end else begin
                                if (6'h2b == _T_263) begin
                                  mem_43 <= _GEN_22;
                                end else begin
                                  if (6'h2b == _T_258) begin
                                    mem_43 <= _GEN_21;
                                  end else begin
                                    if (6'h2b == _T_253) begin
                                      mem_43 <= _GEN_20;
                                    end else begin
                                      if (6'h2b == _T_248) begin
                                        mem_43 <= _GEN_19;
                                      end else begin
                                        if (6'h2b == _T_243) begin
                                          mem_43 <= _GEN_18;
                                        end else begin
                                          if (6'h2b == _T_238) begin
                                            mem_43 <= _GEN_17;
                                          end else begin
                                            if (6'h2b == _T_233) begin
                                              mem_43 <= _GEN_16;
                                            end else begin
                                              if (6'h2b == _T_228) begin
                                                mem_43 <= _GEN_15;
                                              end else begin
                                                if (6'h2b == _T_223) begin
                                                  mem_43 <= _GEN_14;
                                                end else begin
                                                  if (6'h2b == _T_218) begin
                                                    mem_43 <= _GEN_13;
                                                  end else begin
                                                    if (6'h2b == _T_213) begin
                                                      mem_43 <= _GEN_12;
                                                    end else begin
                                                      if (6'h2b == _T_208) begin
                                                        mem_43 <= _GEN_11;
                                                      end else begin
                                                        if (6'h2b == _T_203) begin
                                                          mem_43 <= _GEN_10;
                                                        end else begin
                                                          if (6'h2b == _T_198) begin
                                                            mem_43 <= _GEN_9;
                                                          end else begin
                                                            if (6'h2b == _T_193) begin
                                                              mem_43 <= _GEN_8;
                                                            end else begin
                                                              if (6'h2b == _T_188) begin
                                                                mem_43 <= _GEN_7;
                                                              end else begin
                                                                if (6'h2b == _T_183) begin
                                                                  mem_43 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h2b == _T_178) begin
                                                                    mem_43 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h2b == _T_173) begin
                                                                      mem_43 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h2b == _T_168) begin
                                                                        mem_43 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h2b == _T_163) begin
                                                                          mem_43 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h2b == _T_158) begin
                                                                            mem_43 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h2b == _T_153) begin
                                                                              mem_43 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h2b == _T_308) begin
              mem_43 <= _GEN_31;
            end else begin
              if (6'h2b == _T_303) begin
                mem_43 <= _GEN_30;
              end else begin
                if (6'h2b == _T_298) begin
                  mem_43 <= _GEN_29;
                end else begin
                  if (6'h2b == _T_293) begin
                    mem_43 <= _GEN_28;
                  end else begin
                    if (6'h2b == _T_288) begin
                      mem_43 <= _GEN_27;
                    end else begin
                      if (6'h2b == _T_283) begin
                        mem_43 <= _GEN_26;
                      end else begin
                        if (6'h2b == _T_278) begin
                          mem_43 <= _GEN_25;
                        end else begin
                          if (6'h2b == _T_273) begin
                            mem_43 <= _GEN_24;
                          end else begin
                            if (6'h2b == _T_268) begin
                              mem_43 <= _GEN_23;
                            end else begin
                              if (6'h2b == _T_263) begin
                                mem_43 <= _GEN_22;
                              end else begin
                                if (6'h2b == _T_258) begin
                                  mem_43 <= _GEN_21;
                                end else begin
                                  if (6'h2b == _T_253) begin
                                    mem_43 <= _GEN_20;
                                  end else begin
                                    if (6'h2b == _T_248) begin
                                      mem_43 <= _GEN_19;
                                    end else begin
                                      if (6'h2b == _T_243) begin
                                        mem_43 <= _GEN_18;
                                      end else begin
                                        if (6'h2b == _T_238) begin
                                          mem_43 <= _GEN_17;
                                        end else begin
                                          if (6'h2b == _T_233) begin
                                            mem_43 <= _GEN_16;
                                          end else begin
                                            if (6'h2b == _T_228) begin
                                              mem_43 <= _GEN_15;
                                            end else begin
                                              if (6'h2b == _T_223) begin
                                                mem_43 <= _GEN_14;
                                              end else begin
                                                if (6'h2b == _T_218) begin
                                                  mem_43 <= _GEN_13;
                                                end else begin
                                                  if (6'h2b == _T_213) begin
                                                    mem_43 <= _GEN_12;
                                                  end else begin
                                                    if (6'h2b == _T_208) begin
                                                      mem_43 <= _GEN_11;
                                                    end else begin
                                                      if (6'h2b == _T_203) begin
                                                        mem_43 <= _GEN_10;
                                                      end else begin
                                                        if (6'h2b == _T_198) begin
                                                          mem_43 <= _GEN_9;
                                                        end else begin
                                                          if (6'h2b == _T_193) begin
                                                            mem_43 <= _GEN_8;
                                                          end else begin
                                                            if (6'h2b == _T_188) begin
                                                              mem_43 <= _GEN_7;
                                                            end else begin
                                                              if (6'h2b == _T_183) begin
                                                                mem_43 <= _GEN_6;
                                                              end else begin
                                                                if (6'h2b == _T_178) begin
                                                                  mem_43 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h2b == _T_173) begin
                                                                    mem_43 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h2b == _T_168) begin
                                                                      mem_43 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h2b == _T_163) begin
                                                                        mem_43 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h2b == _T_158) begin
                                                                          mem_43 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h2b == _T_153) begin
                                                                            mem_43 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h2b == _T_308) begin
            mem_43 <= _GEN_31;
          end else begin
            if (6'h2b == _T_303) begin
              mem_43 <= _GEN_30;
            end else begin
              if (6'h2b == _T_298) begin
                mem_43 <= _GEN_29;
              end else begin
                if (6'h2b == _T_293) begin
                  mem_43 <= _GEN_28;
                end else begin
                  if (6'h2b == _T_288) begin
                    mem_43 <= _GEN_27;
                  end else begin
                    if (6'h2b == _T_283) begin
                      mem_43 <= _GEN_26;
                    end else begin
                      if (6'h2b == _T_278) begin
                        mem_43 <= _GEN_25;
                      end else begin
                        if (6'h2b == _T_273) begin
                          mem_43 <= _GEN_24;
                        end else begin
                          if (6'h2b == _T_268) begin
                            mem_43 <= _GEN_23;
                          end else begin
                            if (6'h2b == _T_263) begin
                              mem_43 <= _GEN_22;
                            end else begin
                              if (6'h2b == _T_258) begin
                                mem_43 <= _GEN_21;
                              end else begin
                                if (6'h2b == _T_253) begin
                                  mem_43 <= _GEN_20;
                                end else begin
                                  if (6'h2b == _T_248) begin
                                    mem_43 <= _GEN_19;
                                  end else begin
                                    if (6'h2b == _T_243) begin
                                      mem_43 <= _GEN_18;
                                    end else begin
                                      if (6'h2b == _T_238) begin
                                        mem_43 <= _GEN_17;
                                      end else begin
                                        if (6'h2b == _T_233) begin
                                          mem_43 <= _GEN_16;
                                        end else begin
                                          if (6'h2b == _T_228) begin
                                            mem_43 <= _GEN_15;
                                          end else begin
                                            if (6'h2b == _T_223) begin
                                              mem_43 <= _GEN_14;
                                            end else begin
                                              if (6'h2b == _T_218) begin
                                                mem_43 <= _GEN_13;
                                              end else begin
                                                if (6'h2b == _T_213) begin
                                                  mem_43 <= _GEN_12;
                                                end else begin
                                                  if (6'h2b == _T_208) begin
                                                    mem_43 <= _GEN_11;
                                                  end else begin
                                                    if (6'h2b == _T_203) begin
                                                      mem_43 <= _GEN_10;
                                                    end else begin
                                                      if (6'h2b == _T_198) begin
                                                        mem_43 <= _GEN_9;
                                                      end else begin
                                                        if (6'h2b == _T_193) begin
                                                          mem_43 <= _GEN_8;
                                                        end else begin
                                                          if (6'h2b == _T_188) begin
                                                            mem_43 <= _GEN_7;
                                                          end else begin
                                                            if (6'h2b == _T_183) begin
                                                              mem_43 <= _GEN_6;
                                                            end else begin
                                                              if (6'h2b == _T_178) begin
                                                                mem_43 <= _GEN_5;
                                                              end else begin
                                                                if (6'h2b == _T_173) begin
                                                                  mem_43 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h2b == _T_168) begin
                                                                    mem_43 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h2b == _T_163) begin
                                                                      mem_43 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h2b == _T_158) begin
                                                                        mem_43 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h2b == _T_153) begin
                                                                          mem_43 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h2b == _T_308) begin
          mem_43 <= _GEN_31;
        end else begin
          if (6'h2b == _T_303) begin
            mem_43 <= _GEN_30;
          end else begin
            if (6'h2b == _T_298) begin
              mem_43 <= _GEN_29;
            end else begin
              if (6'h2b == _T_293) begin
                mem_43 <= _GEN_28;
              end else begin
                if (6'h2b == _T_288) begin
                  mem_43 <= _GEN_27;
                end else begin
                  if (6'h2b == _T_283) begin
                    mem_43 <= _GEN_26;
                  end else begin
                    if (6'h2b == _T_278) begin
                      mem_43 <= _GEN_25;
                    end else begin
                      if (6'h2b == _T_273) begin
                        mem_43 <= _GEN_24;
                      end else begin
                        if (6'h2b == _T_268) begin
                          mem_43 <= _GEN_23;
                        end else begin
                          if (6'h2b == _T_263) begin
                            mem_43 <= _GEN_22;
                          end else begin
                            if (6'h2b == _T_258) begin
                              mem_43 <= _GEN_21;
                            end else begin
                              if (6'h2b == _T_253) begin
                                mem_43 <= _GEN_20;
                              end else begin
                                if (6'h2b == _T_248) begin
                                  mem_43 <= _GEN_19;
                                end else begin
                                  if (6'h2b == _T_243) begin
                                    mem_43 <= _GEN_18;
                                  end else begin
                                    if (6'h2b == _T_238) begin
                                      mem_43 <= _GEN_17;
                                    end else begin
                                      if (6'h2b == _T_233) begin
                                        mem_43 <= _GEN_16;
                                      end else begin
                                        if (6'h2b == _T_228) begin
                                          mem_43 <= _GEN_15;
                                        end else begin
                                          if (6'h2b == _T_223) begin
                                            mem_43 <= _GEN_14;
                                          end else begin
                                            if (6'h2b == _T_218) begin
                                              mem_43 <= _GEN_13;
                                            end else begin
                                              if (6'h2b == _T_213) begin
                                                mem_43 <= _GEN_12;
                                              end else begin
                                                if (6'h2b == _T_208) begin
                                                  mem_43 <= _GEN_11;
                                                end else begin
                                                  if (6'h2b == _T_203) begin
                                                    mem_43 <= _GEN_10;
                                                  end else begin
                                                    if (6'h2b == _T_198) begin
                                                      mem_43 <= _GEN_9;
                                                    end else begin
                                                      if (6'h2b == _T_193) begin
                                                        mem_43 <= _GEN_8;
                                                      end else begin
                                                        if (6'h2b == _T_188) begin
                                                          mem_43 <= _GEN_7;
                                                        end else begin
                                                          if (6'h2b == _T_183) begin
                                                            mem_43 <= _GEN_6;
                                                          end else begin
                                                            if (6'h2b == _T_178) begin
                                                              mem_43 <= _GEN_5;
                                                            end else begin
                                                              if (6'h2b == _T_173) begin
                                                                mem_43 <= _GEN_4;
                                                              end else begin
                                                                if (6'h2b == _T_168) begin
                                                                  mem_43 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h2b == _T_163) begin
                                                                    mem_43 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h2b == _T_158) begin
                                                                      mem_43 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h2b == _T_153) begin
                                                                        mem_43 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h2c == wPos) begin
            mem_44 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h2c == _T_308) begin
                mem_44 <= _GEN_31;
              end else begin
                if (6'h2c == _T_303) begin
                  mem_44 <= _GEN_30;
                end else begin
                  if (6'h2c == _T_298) begin
                    mem_44 <= _GEN_29;
                  end else begin
                    if (6'h2c == _T_293) begin
                      mem_44 <= _GEN_28;
                    end else begin
                      if (6'h2c == _T_288) begin
                        mem_44 <= _GEN_27;
                      end else begin
                        if (6'h2c == _T_283) begin
                          mem_44 <= _GEN_26;
                        end else begin
                          if (6'h2c == _T_278) begin
                            mem_44 <= _GEN_25;
                          end else begin
                            if (6'h2c == _T_273) begin
                              mem_44 <= _GEN_24;
                            end else begin
                              if (6'h2c == _T_268) begin
                                mem_44 <= _GEN_23;
                              end else begin
                                if (6'h2c == _T_263) begin
                                  mem_44 <= _GEN_22;
                                end else begin
                                  if (6'h2c == _T_258) begin
                                    mem_44 <= _GEN_21;
                                  end else begin
                                    if (6'h2c == _T_253) begin
                                      mem_44 <= _GEN_20;
                                    end else begin
                                      if (6'h2c == _T_248) begin
                                        mem_44 <= _GEN_19;
                                      end else begin
                                        if (6'h2c == _T_243) begin
                                          mem_44 <= _GEN_18;
                                        end else begin
                                          if (6'h2c == _T_238) begin
                                            mem_44 <= _GEN_17;
                                          end else begin
                                            if (6'h2c == _T_233) begin
                                              mem_44 <= _GEN_16;
                                            end else begin
                                              if (6'h2c == _T_228) begin
                                                mem_44 <= _GEN_15;
                                              end else begin
                                                if (6'h2c == _T_223) begin
                                                  mem_44 <= _GEN_14;
                                                end else begin
                                                  if (6'h2c == _T_218) begin
                                                    mem_44 <= _GEN_13;
                                                  end else begin
                                                    if (6'h2c == _T_213) begin
                                                      mem_44 <= _GEN_12;
                                                    end else begin
                                                      if (6'h2c == _T_208) begin
                                                        mem_44 <= _GEN_11;
                                                      end else begin
                                                        if (6'h2c == _T_203) begin
                                                          mem_44 <= _GEN_10;
                                                        end else begin
                                                          if (6'h2c == _T_198) begin
                                                            mem_44 <= _GEN_9;
                                                          end else begin
                                                            if (6'h2c == _T_193) begin
                                                              mem_44 <= _GEN_8;
                                                            end else begin
                                                              if (6'h2c == _T_188) begin
                                                                mem_44 <= _GEN_7;
                                                              end else begin
                                                                if (6'h2c == _T_183) begin
                                                                  mem_44 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h2c == _T_178) begin
                                                                    mem_44 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h2c == _T_173) begin
                                                                      mem_44 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h2c == _T_168) begin
                                                                        mem_44 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h2c == _T_163) begin
                                                                          mem_44 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h2c == _T_158) begin
                                                                            mem_44 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h2c == _T_153) begin
                                                                              mem_44 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h2c == _T_308) begin
              mem_44 <= _GEN_31;
            end else begin
              if (6'h2c == _T_303) begin
                mem_44 <= _GEN_30;
              end else begin
                if (6'h2c == _T_298) begin
                  mem_44 <= _GEN_29;
                end else begin
                  if (6'h2c == _T_293) begin
                    mem_44 <= _GEN_28;
                  end else begin
                    if (6'h2c == _T_288) begin
                      mem_44 <= _GEN_27;
                    end else begin
                      if (6'h2c == _T_283) begin
                        mem_44 <= _GEN_26;
                      end else begin
                        if (6'h2c == _T_278) begin
                          mem_44 <= _GEN_25;
                        end else begin
                          if (6'h2c == _T_273) begin
                            mem_44 <= _GEN_24;
                          end else begin
                            if (6'h2c == _T_268) begin
                              mem_44 <= _GEN_23;
                            end else begin
                              if (6'h2c == _T_263) begin
                                mem_44 <= _GEN_22;
                              end else begin
                                if (6'h2c == _T_258) begin
                                  mem_44 <= _GEN_21;
                                end else begin
                                  if (6'h2c == _T_253) begin
                                    mem_44 <= _GEN_20;
                                  end else begin
                                    if (6'h2c == _T_248) begin
                                      mem_44 <= _GEN_19;
                                    end else begin
                                      if (6'h2c == _T_243) begin
                                        mem_44 <= _GEN_18;
                                      end else begin
                                        if (6'h2c == _T_238) begin
                                          mem_44 <= _GEN_17;
                                        end else begin
                                          if (6'h2c == _T_233) begin
                                            mem_44 <= _GEN_16;
                                          end else begin
                                            if (6'h2c == _T_228) begin
                                              mem_44 <= _GEN_15;
                                            end else begin
                                              if (6'h2c == _T_223) begin
                                                mem_44 <= _GEN_14;
                                              end else begin
                                                if (6'h2c == _T_218) begin
                                                  mem_44 <= _GEN_13;
                                                end else begin
                                                  if (6'h2c == _T_213) begin
                                                    mem_44 <= _GEN_12;
                                                  end else begin
                                                    if (6'h2c == _T_208) begin
                                                      mem_44 <= _GEN_11;
                                                    end else begin
                                                      if (6'h2c == _T_203) begin
                                                        mem_44 <= _GEN_10;
                                                      end else begin
                                                        if (6'h2c == _T_198) begin
                                                          mem_44 <= _GEN_9;
                                                        end else begin
                                                          if (6'h2c == _T_193) begin
                                                            mem_44 <= _GEN_8;
                                                          end else begin
                                                            if (6'h2c == _T_188) begin
                                                              mem_44 <= _GEN_7;
                                                            end else begin
                                                              if (6'h2c == _T_183) begin
                                                                mem_44 <= _GEN_6;
                                                              end else begin
                                                                if (6'h2c == _T_178) begin
                                                                  mem_44 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h2c == _T_173) begin
                                                                    mem_44 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h2c == _T_168) begin
                                                                      mem_44 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h2c == _T_163) begin
                                                                        mem_44 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h2c == _T_158) begin
                                                                          mem_44 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h2c == _T_153) begin
                                                                            mem_44 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h2c == _T_308) begin
            mem_44 <= _GEN_31;
          end else begin
            if (6'h2c == _T_303) begin
              mem_44 <= _GEN_30;
            end else begin
              if (6'h2c == _T_298) begin
                mem_44 <= _GEN_29;
              end else begin
                if (6'h2c == _T_293) begin
                  mem_44 <= _GEN_28;
                end else begin
                  if (6'h2c == _T_288) begin
                    mem_44 <= _GEN_27;
                  end else begin
                    if (6'h2c == _T_283) begin
                      mem_44 <= _GEN_26;
                    end else begin
                      if (6'h2c == _T_278) begin
                        mem_44 <= _GEN_25;
                      end else begin
                        if (6'h2c == _T_273) begin
                          mem_44 <= _GEN_24;
                        end else begin
                          if (6'h2c == _T_268) begin
                            mem_44 <= _GEN_23;
                          end else begin
                            if (6'h2c == _T_263) begin
                              mem_44 <= _GEN_22;
                            end else begin
                              if (6'h2c == _T_258) begin
                                mem_44 <= _GEN_21;
                              end else begin
                                if (6'h2c == _T_253) begin
                                  mem_44 <= _GEN_20;
                                end else begin
                                  if (6'h2c == _T_248) begin
                                    mem_44 <= _GEN_19;
                                  end else begin
                                    if (6'h2c == _T_243) begin
                                      mem_44 <= _GEN_18;
                                    end else begin
                                      if (6'h2c == _T_238) begin
                                        mem_44 <= _GEN_17;
                                      end else begin
                                        if (6'h2c == _T_233) begin
                                          mem_44 <= _GEN_16;
                                        end else begin
                                          if (6'h2c == _T_228) begin
                                            mem_44 <= _GEN_15;
                                          end else begin
                                            if (6'h2c == _T_223) begin
                                              mem_44 <= _GEN_14;
                                            end else begin
                                              if (6'h2c == _T_218) begin
                                                mem_44 <= _GEN_13;
                                              end else begin
                                                if (6'h2c == _T_213) begin
                                                  mem_44 <= _GEN_12;
                                                end else begin
                                                  if (6'h2c == _T_208) begin
                                                    mem_44 <= _GEN_11;
                                                  end else begin
                                                    if (6'h2c == _T_203) begin
                                                      mem_44 <= _GEN_10;
                                                    end else begin
                                                      if (6'h2c == _T_198) begin
                                                        mem_44 <= _GEN_9;
                                                      end else begin
                                                        if (6'h2c == _T_193) begin
                                                          mem_44 <= _GEN_8;
                                                        end else begin
                                                          if (6'h2c == _T_188) begin
                                                            mem_44 <= _GEN_7;
                                                          end else begin
                                                            if (6'h2c == _T_183) begin
                                                              mem_44 <= _GEN_6;
                                                            end else begin
                                                              if (6'h2c == _T_178) begin
                                                                mem_44 <= _GEN_5;
                                                              end else begin
                                                                if (6'h2c == _T_173) begin
                                                                  mem_44 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h2c == _T_168) begin
                                                                    mem_44 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h2c == _T_163) begin
                                                                      mem_44 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h2c == _T_158) begin
                                                                        mem_44 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h2c == _T_153) begin
                                                                          mem_44 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h2c == _T_308) begin
          mem_44 <= _GEN_31;
        end else begin
          if (6'h2c == _T_303) begin
            mem_44 <= _GEN_30;
          end else begin
            if (6'h2c == _T_298) begin
              mem_44 <= _GEN_29;
            end else begin
              if (6'h2c == _T_293) begin
                mem_44 <= _GEN_28;
              end else begin
                if (6'h2c == _T_288) begin
                  mem_44 <= _GEN_27;
                end else begin
                  if (6'h2c == _T_283) begin
                    mem_44 <= _GEN_26;
                  end else begin
                    if (6'h2c == _T_278) begin
                      mem_44 <= _GEN_25;
                    end else begin
                      if (6'h2c == _T_273) begin
                        mem_44 <= _GEN_24;
                      end else begin
                        if (6'h2c == _T_268) begin
                          mem_44 <= _GEN_23;
                        end else begin
                          if (6'h2c == _T_263) begin
                            mem_44 <= _GEN_22;
                          end else begin
                            if (6'h2c == _T_258) begin
                              mem_44 <= _GEN_21;
                            end else begin
                              if (6'h2c == _T_253) begin
                                mem_44 <= _GEN_20;
                              end else begin
                                if (6'h2c == _T_248) begin
                                  mem_44 <= _GEN_19;
                                end else begin
                                  if (6'h2c == _T_243) begin
                                    mem_44 <= _GEN_18;
                                  end else begin
                                    if (6'h2c == _T_238) begin
                                      mem_44 <= _GEN_17;
                                    end else begin
                                      if (6'h2c == _T_233) begin
                                        mem_44 <= _GEN_16;
                                      end else begin
                                        if (6'h2c == _T_228) begin
                                          mem_44 <= _GEN_15;
                                        end else begin
                                          if (6'h2c == _T_223) begin
                                            mem_44 <= _GEN_14;
                                          end else begin
                                            if (6'h2c == _T_218) begin
                                              mem_44 <= _GEN_13;
                                            end else begin
                                              if (6'h2c == _T_213) begin
                                                mem_44 <= _GEN_12;
                                              end else begin
                                                if (6'h2c == _T_208) begin
                                                  mem_44 <= _GEN_11;
                                                end else begin
                                                  if (6'h2c == _T_203) begin
                                                    mem_44 <= _GEN_10;
                                                  end else begin
                                                    if (6'h2c == _T_198) begin
                                                      mem_44 <= _GEN_9;
                                                    end else begin
                                                      if (6'h2c == _T_193) begin
                                                        mem_44 <= _GEN_8;
                                                      end else begin
                                                        if (6'h2c == _T_188) begin
                                                          mem_44 <= _GEN_7;
                                                        end else begin
                                                          if (6'h2c == _T_183) begin
                                                            mem_44 <= _GEN_6;
                                                          end else begin
                                                            if (6'h2c == _T_178) begin
                                                              mem_44 <= _GEN_5;
                                                            end else begin
                                                              if (6'h2c == _T_173) begin
                                                                mem_44 <= _GEN_4;
                                                              end else begin
                                                                if (6'h2c == _T_168) begin
                                                                  mem_44 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h2c == _T_163) begin
                                                                    mem_44 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h2c == _T_158) begin
                                                                      mem_44 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h2c == _T_153) begin
                                                                        mem_44 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h2d == wPos) begin
            mem_45 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h2d == _T_308) begin
                mem_45 <= _GEN_31;
              end else begin
                if (6'h2d == _T_303) begin
                  mem_45 <= _GEN_30;
                end else begin
                  if (6'h2d == _T_298) begin
                    mem_45 <= _GEN_29;
                  end else begin
                    if (6'h2d == _T_293) begin
                      mem_45 <= _GEN_28;
                    end else begin
                      if (6'h2d == _T_288) begin
                        mem_45 <= _GEN_27;
                      end else begin
                        if (6'h2d == _T_283) begin
                          mem_45 <= _GEN_26;
                        end else begin
                          if (6'h2d == _T_278) begin
                            mem_45 <= _GEN_25;
                          end else begin
                            if (6'h2d == _T_273) begin
                              mem_45 <= _GEN_24;
                            end else begin
                              if (6'h2d == _T_268) begin
                                mem_45 <= _GEN_23;
                              end else begin
                                if (6'h2d == _T_263) begin
                                  mem_45 <= _GEN_22;
                                end else begin
                                  if (6'h2d == _T_258) begin
                                    mem_45 <= _GEN_21;
                                  end else begin
                                    if (6'h2d == _T_253) begin
                                      mem_45 <= _GEN_20;
                                    end else begin
                                      if (6'h2d == _T_248) begin
                                        mem_45 <= _GEN_19;
                                      end else begin
                                        if (6'h2d == _T_243) begin
                                          mem_45 <= _GEN_18;
                                        end else begin
                                          if (6'h2d == _T_238) begin
                                            mem_45 <= _GEN_17;
                                          end else begin
                                            if (6'h2d == _T_233) begin
                                              mem_45 <= _GEN_16;
                                            end else begin
                                              if (6'h2d == _T_228) begin
                                                mem_45 <= _GEN_15;
                                              end else begin
                                                if (6'h2d == _T_223) begin
                                                  mem_45 <= _GEN_14;
                                                end else begin
                                                  if (6'h2d == _T_218) begin
                                                    mem_45 <= _GEN_13;
                                                  end else begin
                                                    if (6'h2d == _T_213) begin
                                                      mem_45 <= _GEN_12;
                                                    end else begin
                                                      if (6'h2d == _T_208) begin
                                                        mem_45 <= _GEN_11;
                                                      end else begin
                                                        if (6'h2d == _T_203) begin
                                                          mem_45 <= _GEN_10;
                                                        end else begin
                                                          if (6'h2d == _T_198) begin
                                                            mem_45 <= _GEN_9;
                                                          end else begin
                                                            if (6'h2d == _T_193) begin
                                                              mem_45 <= _GEN_8;
                                                            end else begin
                                                              if (6'h2d == _T_188) begin
                                                                mem_45 <= _GEN_7;
                                                              end else begin
                                                                if (6'h2d == _T_183) begin
                                                                  mem_45 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h2d == _T_178) begin
                                                                    mem_45 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h2d == _T_173) begin
                                                                      mem_45 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h2d == _T_168) begin
                                                                        mem_45 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h2d == _T_163) begin
                                                                          mem_45 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h2d == _T_158) begin
                                                                            mem_45 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h2d == _T_153) begin
                                                                              mem_45 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h2d == _T_308) begin
              mem_45 <= _GEN_31;
            end else begin
              if (6'h2d == _T_303) begin
                mem_45 <= _GEN_30;
              end else begin
                if (6'h2d == _T_298) begin
                  mem_45 <= _GEN_29;
                end else begin
                  if (6'h2d == _T_293) begin
                    mem_45 <= _GEN_28;
                  end else begin
                    if (6'h2d == _T_288) begin
                      mem_45 <= _GEN_27;
                    end else begin
                      if (6'h2d == _T_283) begin
                        mem_45 <= _GEN_26;
                      end else begin
                        if (6'h2d == _T_278) begin
                          mem_45 <= _GEN_25;
                        end else begin
                          if (6'h2d == _T_273) begin
                            mem_45 <= _GEN_24;
                          end else begin
                            if (6'h2d == _T_268) begin
                              mem_45 <= _GEN_23;
                            end else begin
                              if (6'h2d == _T_263) begin
                                mem_45 <= _GEN_22;
                              end else begin
                                if (6'h2d == _T_258) begin
                                  mem_45 <= _GEN_21;
                                end else begin
                                  if (6'h2d == _T_253) begin
                                    mem_45 <= _GEN_20;
                                  end else begin
                                    if (6'h2d == _T_248) begin
                                      mem_45 <= _GEN_19;
                                    end else begin
                                      if (6'h2d == _T_243) begin
                                        mem_45 <= _GEN_18;
                                      end else begin
                                        if (6'h2d == _T_238) begin
                                          mem_45 <= _GEN_17;
                                        end else begin
                                          if (6'h2d == _T_233) begin
                                            mem_45 <= _GEN_16;
                                          end else begin
                                            if (6'h2d == _T_228) begin
                                              mem_45 <= _GEN_15;
                                            end else begin
                                              if (6'h2d == _T_223) begin
                                                mem_45 <= _GEN_14;
                                              end else begin
                                                if (6'h2d == _T_218) begin
                                                  mem_45 <= _GEN_13;
                                                end else begin
                                                  if (6'h2d == _T_213) begin
                                                    mem_45 <= _GEN_12;
                                                  end else begin
                                                    if (6'h2d == _T_208) begin
                                                      mem_45 <= _GEN_11;
                                                    end else begin
                                                      if (6'h2d == _T_203) begin
                                                        mem_45 <= _GEN_10;
                                                      end else begin
                                                        if (6'h2d == _T_198) begin
                                                          mem_45 <= _GEN_9;
                                                        end else begin
                                                          if (6'h2d == _T_193) begin
                                                            mem_45 <= _GEN_8;
                                                          end else begin
                                                            if (6'h2d == _T_188) begin
                                                              mem_45 <= _GEN_7;
                                                            end else begin
                                                              if (6'h2d == _T_183) begin
                                                                mem_45 <= _GEN_6;
                                                              end else begin
                                                                if (6'h2d == _T_178) begin
                                                                  mem_45 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h2d == _T_173) begin
                                                                    mem_45 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h2d == _T_168) begin
                                                                      mem_45 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h2d == _T_163) begin
                                                                        mem_45 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h2d == _T_158) begin
                                                                          mem_45 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h2d == _T_153) begin
                                                                            mem_45 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h2d == _T_308) begin
            mem_45 <= _GEN_31;
          end else begin
            if (6'h2d == _T_303) begin
              mem_45 <= _GEN_30;
            end else begin
              if (6'h2d == _T_298) begin
                mem_45 <= _GEN_29;
              end else begin
                if (6'h2d == _T_293) begin
                  mem_45 <= _GEN_28;
                end else begin
                  if (6'h2d == _T_288) begin
                    mem_45 <= _GEN_27;
                  end else begin
                    if (6'h2d == _T_283) begin
                      mem_45 <= _GEN_26;
                    end else begin
                      if (6'h2d == _T_278) begin
                        mem_45 <= _GEN_25;
                      end else begin
                        if (6'h2d == _T_273) begin
                          mem_45 <= _GEN_24;
                        end else begin
                          if (6'h2d == _T_268) begin
                            mem_45 <= _GEN_23;
                          end else begin
                            if (6'h2d == _T_263) begin
                              mem_45 <= _GEN_22;
                            end else begin
                              if (6'h2d == _T_258) begin
                                mem_45 <= _GEN_21;
                              end else begin
                                if (6'h2d == _T_253) begin
                                  mem_45 <= _GEN_20;
                                end else begin
                                  if (6'h2d == _T_248) begin
                                    mem_45 <= _GEN_19;
                                  end else begin
                                    if (6'h2d == _T_243) begin
                                      mem_45 <= _GEN_18;
                                    end else begin
                                      if (6'h2d == _T_238) begin
                                        mem_45 <= _GEN_17;
                                      end else begin
                                        if (6'h2d == _T_233) begin
                                          mem_45 <= _GEN_16;
                                        end else begin
                                          if (6'h2d == _T_228) begin
                                            mem_45 <= _GEN_15;
                                          end else begin
                                            if (6'h2d == _T_223) begin
                                              mem_45 <= _GEN_14;
                                            end else begin
                                              if (6'h2d == _T_218) begin
                                                mem_45 <= _GEN_13;
                                              end else begin
                                                if (6'h2d == _T_213) begin
                                                  mem_45 <= _GEN_12;
                                                end else begin
                                                  if (6'h2d == _T_208) begin
                                                    mem_45 <= _GEN_11;
                                                  end else begin
                                                    if (6'h2d == _T_203) begin
                                                      mem_45 <= _GEN_10;
                                                    end else begin
                                                      if (6'h2d == _T_198) begin
                                                        mem_45 <= _GEN_9;
                                                      end else begin
                                                        if (6'h2d == _T_193) begin
                                                          mem_45 <= _GEN_8;
                                                        end else begin
                                                          if (6'h2d == _T_188) begin
                                                            mem_45 <= _GEN_7;
                                                          end else begin
                                                            if (6'h2d == _T_183) begin
                                                              mem_45 <= _GEN_6;
                                                            end else begin
                                                              if (6'h2d == _T_178) begin
                                                                mem_45 <= _GEN_5;
                                                              end else begin
                                                                if (6'h2d == _T_173) begin
                                                                  mem_45 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h2d == _T_168) begin
                                                                    mem_45 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h2d == _T_163) begin
                                                                      mem_45 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h2d == _T_158) begin
                                                                        mem_45 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h2d == _T_153) begin
                                                                          mem_45 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h2d == _T_308) begin
          mem_45 <= _GEN_31;
        end else begin
          if (6'h2d == _T_303) begin
            mem_45 <= _GEN_30;
          end else begin
            if (6'h2d == _T_298) begin
              mem_45 <= _GEN_29;
            end else begin
              if (6'h2d == _T_293) begin
                mem_45 <= _GEN_28;
              end else begin
                if (6'h2d == _T_288) begin
                  mem_45 <= _GEN_27;
                end else begin
                  if (6'h2d == _T_283) begin
                    mem_45 <= _GEN_26;
                  end else begin
                    if (6'h2d == _T_278) begin
                      mem_45 <= _GEN_25;
                    end else begin
                      if (6'h2d == _T_273) begin
                        mem_45 <= _GEN_24;
                      end else begin
                        if (6'h2d == _T_268) begin
                          mem_45 <= _GEN_23;
                        end else begin
                          if (6'h2d == _T_263) begin
                            mem_45 <= _GEN_22;
                          end else begin
                            if (6'h2d == _T_258) begin
                              mem_45 <= _GEN_21;
                            end else begin
                              if (6'h2d == _T_253) begin
                                mem_45 <= _GEN_20;
                              end else begin
                                if (6'h2d == _T_248) begin
                                  mem_45 <= _GEN_19;
                                end else begin
                                  if (6'h2d == _T_243) begin
                                    mem_45 <= _GEN_18;
                                  end else begin
                                    if (6'h2d == _T_238) begin
                                      mem_45 <= _GEN_17;
                                    end else begin
                                      if (6'h2d == _T_233) begin
                                        mem_45 <= _GEN_16;
                                      end else begin
                                        if (6'h2d == _T_228) begin
                                          mem_45 <= _GEN_15;
                                        end else begin
                                          if (6'h2d == _T_223) begin
                                            mem_45 <= _GEN_14;
                                          end else begin
                                            if (6'h2d == _T_218) begin
                                              mem_45 <= _GEN_13;
                                            end else begin
                                              if (6'h2d == _T_213) begin
                                                mem_45 <= _GEN_12;
                                              end else begin
                                                if (6'h2d == _T_208) begin
                                                  mem_45 <= _GEN_11;
                                                end else begin
                                                  if (6'h2d == _T_203) begin
                                                    mem_45 <= _GEN_10;
                                                  end else begin
                                                    if (6'h2d == _T_198) begin
                                                      mem_45 <= _GEN_9;
                                                    end else begin
                                                      if (6'h2d == _T_193) begin
                                                        mem_45 <= _GEN_8;
                                                      end else begin
                                                        if (6'h2d == _T_188) begin
                                                          mem_45 <= _GEN_7;
                                                        end else begin
                                                          if (6'h2d == _T_183) begin
                                                            mem_45 <= _GEN_6;
                                                          end else begin
                                                            if (6'h2d == _T_178) begin
                                                              mem_45 <= _GEN_5;
                                                            end else begin
                                                              if (6'h2d == _T_173) begin
                                                                mem_45 <= _GEN_4;
                                                              end else begin
                                                                if (6'h2d == _T_168) begin
                                                                  mem_45 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h2d == _T_163) begin
                                                                    mem_45 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h2d == _T_158) begin
                                                                      mem_45 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h2d == _T_153) begin
                                                                        mem_45 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h2e == wPos) begin
            mem_46 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h2e == _T_308) begin
                mem_46 <= _GEN_31;
              end else begin
                if (6'h2e == _T_303) begin
                  mem_46 <= _GEN_30;
                end else begin
                  if (6'h2e == _T_298) begin
                    mem_46 <= _GEN_29;
                  end else begin
                    if (6'h2e == _T_293) begin
                      mem_46 <= _GEN_28;
                    end else begin
                      if (6'h2e == _T_288) begin
                        mem_46 <= _GEN_27;
                      end else begin
                        if (6'h2e == _T_283) begin
                          mem_46 <= _GEN_26;
                        end else begin
                          if (6'h2e == _T_278) begin
                            mem_46 <= _GEN_25;
                          end else begin
                            if (6'h2e == _T_273) begin
                              mem_46 <= _GEN_24;
                            end else begin
                              if (6'h2e == _T_268) begin
                                mem_46 <= _GEN_23;
                              end else begin
                                if (6'h2e == _T_263) begin
                                  mem_46 <= _GEN_22;
                                end else begin
                                  if (6'h2e == _T_258) begin
                                    mem_46 <= _GEN_21;
                                  end else begin
                                    if (6'h2e == _T_253) begin
                                      mem_46 <= _GEN_20;
                                    end else begin
                                      if (6'h2e == _T_248) begin
                                        mem_46 <= _GEN_19;
                                      end else begin
                                        if (6'h2e == _T_243) begin
                                          mem_46 <= _GEN_18;
                                        end else begin
                                          if (6'h2e == _T_238) begin
                                            mem_46 <= _GEN_17;
                                          end else begin
                                            if (6'h2e == _T_233) begin
                                              mem_46 <= _GEN_16;
                                            end else begin
                                              if (6'h2e == _T_228) begin
                                                mem_46 <= _GEN_15;
                                              end else begin
                                                if (6'h2e == _T_223) begin
                                                  mem_46 <= _GEN_14;
                                                end else begin
                                                  if (6'h2e == _T_218) begin
                                                    mem_46 <= _GEN_13;
                                                  end else begin
                                                    if (6'h2e == _T_213) begin
                                                      mem_46 <= _GEN_12;
                                                    end else begin
                                                      if (6'h2e == _T_208) begin
                                                        mem_46 <= _GEN_11;
                                                      end else begin
                                                        if (6'h2e == _T_203) begin
                                                          mem_46 <= _GEN_10;
                                                        end else begin
                                                          if (6'h2e == _T_198) begin
                                                            mem_46 <= _GEN_9;
                                                          end else begin
                                                            if (6'h2e == _T_193) begin
                                                              mem_46 <= _GEN_8;
                                                            end else begin
                                                              if (6'h2e == _T_188) begin
                                                                mem_46 <= _GEN_7;
                                                              end else begin
                                                                if (6'h2e == _T_183) begin
                                                                  mem_46 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h2e == _T_178) begin
                                                                    mem_46 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h2e == _T_173) begin
                                                                      mem_46 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h2e == _T_168) begin
                                                                        mem_46 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h2e == _T_163) begin
                                                                          mem_46 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h2e == _T_158) begin
                                                                            mem_46 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h2e == _T_153) begin
                                                                              mem_46 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h2e == _T_308) begin
              mem_46 <= _GEN_31;
            end else begin
              if (6'h2e == _T_303) begin
                mem_46 <= _GEN_30;
              end else begin
                if (6'h2e == _T_298) begin
                  mem_46 <= _GEN_29;
                end else begin
                  if (6'h2e == _T_293) begin
                    mem_46 <= _GEN_28;
                  end else begin
                    if (6'h2e == _T_288) begin
                      mem_46 <= _GEN_27;
                    end else begin
                      if (6'h2e == _T_283) begin
                        mem_46 <= _GEN_26;
                      end else begin
                        if (6'h2e == _T_278) begin
                          mem_46 <= _GEN_25;
                        end else begin
                          if (6'h2e == _T_273) begin
                            mem_46 <= _GEN_24;
                          end else begin
                            if (6'h2e == _T_268) begin
                              mem_46 <= _GEN_23;
                            end else begin
                              if (6'h2e == _T_263) begin
                                mem_46 <= _GEN_22;
                              end else begin
                                if (6'h2e == _T_258) begin
                                  mem_46 <= _GEN_21;
                                end else begin
                                  if (6'h2e == _T_253) begin
                                    mem_46 <= _GEN_20;
                                  end else begin
                                    if (6'h2e == _T_248) begin
                                      mem_46 <= _GEN_19;
                                    end else begin
                                      if (6'h2e == _T_243) begin
                                        mem_46 <= _GEN_18;
                                      end else begin
                                        if (6'h2e == _T_238) begin
                                          mem_46 <= _GEN_17;
                                        end else begin
                                          if (6'h2e == _T_233) begin
                                            mem_46 <= _GEN_16;
                                          end else begin
                                            if (6'h2e == _T_228) begin
                                              mem_46 <= _GEN_15;
                                            end else begin
                                              if (6'h2e == _T_223) begin
                                                mem_46 <= _GEN_14;
                                              end else begin
                                                if (6'h2e == _T_218) begin
                                                  mem_46 <= _GEN_13;
                                                end else begin
                                                  if (6'h2e == _T_213) begin
                                                    mem_46 <= _GEN_12;
                                                  end else begin
                                                    if (6'h2e == _T_208) begin
                                                      mem_46 <= _GEN_11;
                                                    end else begin
                                                      if (6'h2e == _T_203) begin
                                                        mem_46 <= _GEN_10;
                                                      end else begin
                                                        if (6'h2e == _T_198) begin
                                                          mem_46 <= _GEN_9;
                                                        end else begin
                                                          if (6'h2e == _T_193) begin
                                                            mem_46 <= _GEN_8;
                                                          end else begin
                                                            if (6'h2e == _T_188) begin
                                                              mem_46 <= _GEN_7;
                                                            end else begin
                                                              if (6'h2e == _T_183) begin
                                                                mem_46 <= _GEN_6;
                                                              end else begin
                                                                if (6'h2e == _T_178) begin
                                                                  mem_46 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h2e == _T_173) begin
                                                                    mem_46 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h2e == _T_168) begin
                                                                      mem_46 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h2e == _T_163) begin
                                                                        mem_46 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h2e == _T_158) begin
                                                                          mem_46 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h2e == _T_153) begin
                                                                            mem_46 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h2e == _T_308) begin
            mem_46 <= _GEN_31;
          end else begin
            if (6'h2e == _T_303) begin
              mem_46 <= _GEN_30;
            end else begin
              if (6'h2e == _T_298) begin
                mem_46 <= _GEN_29;
              end else begin
                if (6'h2e == _T_293) begin
                  mem_46 <= _GEN_28;
                end else begin
                  if (6'h2e == _T_288) begin
                    mem_46 <= _GEN_27;
                  end else begin
                    if (6'h2e == _T_283) begin
                      mem_46 <= _GEN_26;
                    end else begin
                      if (6'h2e == _T_278) begin
                        mem_46 <= _GEN_25;
                      end else begin
                        if (6'h2e == _T_273) begin
                          mem_46 <= _GEN_24;
                        end else begin
                          if (6'h2e == _T_268) begin
                            mem_46 <= _GEN_23;
                          end else begin
                            if (6'h2e == _T_263) begin
                              mem_46 <= _GEN_22;
                            end else begin
                              if (6'h2e == _T_258) begin
                                mem_46 <= _GEN_21;
                              end else begin
                                if (6'h2e == _T_253) begin
                                  mem_46 <= _GEN_20;
                                end else begin
                                  if (6'h2e == _T_248) begin
                                    mem_46 <= _GEN_19;
                                  end else begin
                                    if (6'h2e == _T_243) begin
                                      mem_46 <= _GEN_18;
                                    end else begin
                                      if (6'h2e == _T_238) begin
                                        mem_46 <= _GEN_17;
                                      end else begin
                                        if (6'h2e == _T_233) begin
                                          mem_46 <= _GEN_16;
                                        end else begin
                                          if (6'h2e == _T_228) begin
                                            mem_46 <= _GEN_15;
                                          end else begin
                                            if (6'h2e == _T_223) begin
                                              mem_46 <= _GEN_14;
                                            end else begin
                                              if (6'h2e == _T_218) begin
                                                mem_46 <= _GEN_13;
                                              end else begin
                                                if (6'h2e == _T_213) begin
                                                  mem_46 <= _GEN_12;
                                                end else begin
                                                  if (6'h2e == _T_208) begin
                                                    mem_46 <= _GEN_11;
                                                  end else begin
                                                    if (6'h2e == _T_203) begin
                                                      mem_46 <= _GEN_10;
                                                    end else begin
                                                      if (6'h2e == _T_198) begin
                                                        mem_46 <= _GEN_9;
                                                      end else begin
                                                        if (6'h2e == _T_193) begin
                                                          mem_46 <= _GEN_8;
                                                        end else begin
                                                          if (6'h2e == _T_188) begin
                                                            mem_46 <= _GEN_7;
                                                          end else begin
                                                            if (6'h2e == _T_183) begin
                                                              mem_46 <= _GEN_6;
                                                            end else begin
                                                              if (6'h2e == _T_178) begin
                                                                mem_46 <= _GEN_5;
                                                              end else begin
                                                                if (6'h2e == _T_173) begin
                                                                  mem_46 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h2e == _T_168) begin
                                                                    mem_46 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h2e == _T_163) begin
                                                                      mem_46 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h2e == _T_158) begin
                                                                        mem_46 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h2e == _T_153) begin
                                                                          mem_46 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h2e == _T_308) begin
          mem_46 <= _GEN_31;
        end else begin
          if (6'h2e == _T_303) begin
            mem_46 <= _GEN_30;
          end else begin
            if (6'h2e == _T_298) begin
              mem_46 <= _GEN_29;
            end else begin
              if (6'h2e == _T_293) begin
                mem_46 <= _GEN_28;
              end else begin
                if (6'h2e == _T_288) begin
                  mem_46 <= _GEN_27;
                end else begin
                  if (6'h2e == _T_283) begin
                    mem_46 <= _GEN_26;
                  end else begin
                    if (6'h2e == _T_278) begin
                      mem_46 <= _GEN_25;
                    end else begin
                      if (6'h2e == _T_273) begin
                        mem_46 <= _GEN_24;
                      end else begin
                        if (6'h2e == _T_268) begin
                          mem_46 <= _GEN_23;
                        end else begin
                          if (6'h2e == _T_263) begin
                            mem_46 <= _GEN_22;
                          end else begin
                            if (6'h2e == _T_258) begin
                              mem_46 <= _GEN_21;
                            end else begin
                              if (6'h2e == _T_253) begin
                                mem_46 <= _GEN_20;
                              end else begin
                                if (6'h2e == _T_248) begin
                                  mem_46 <= _GEN_19;
                                end else begin
                                  if (6'h2e == _T_243) begin
                                    mem_46 <= _GEN_18;
                                  end else begin
                                    if (6'h2e == _T_238) begin
                                      mem_46 <= _GEN_17;
                                    end else begin
                                      if (6'h2e == _T_233) begin
                                        mem_46 <= _GEN_16;
                                      end else begin
                                        if (6'h2e == _T_228) begin
                                          mem_46 <= _GEN_15;
                                        end else begin
                                          if (6'h2e == _T_223) begin
                                            mem_46 <= _GEN_14;
                                          end else begin
                                            if (6'h2e == _T_218) begin
                                              mem_46 <= _GEN_13;
                                            end else begin
                                              if (6'h2e == _T_213) begin
                                                mem_46 <= _GEN_12;
                                              end else begin
                                                if (6'h2e == _T_208) begin
                                                  mem_46 <= _GEN_11;
                                                end else begin
                                                  if (6'h2e == _T_203) begin
                                                    mem_46 <= _GEN_10;
                                                  end else begin
                                                    if (6'h2e == _T_198) begin
                                                      mem_46 <= _GEN_9;
                                                    end else begin
                                                      if (6'h2e == _T_193) begin
                                                        mem_46 <= _GEN_8;
                                                      end else begin
                                                        if (6'h2e == _T_188) begin
                                                          mem_46 <= _GEN_7;
                                                        end else begin
                                                          if (6'h2e == _T_183) begin
                                                            mem_46 <= _GEN_6;
                                                          end else begin
                                                            if (6'h2e == _T_178) begin
                                                              mem_46 <= _GEN_5;
                                                            end else begin
                                                              if (6'h2e == _T_173) begin
                                                                mem_46 <= _GEN_4;
                                                              end else begin
                                                                if (6'h2e == _T_168) begin
                                                                  mem_46 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h2e == _T_163) begin
                                                                    mem_46 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h2e == _T_158) begin
                                                                      mem_46 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h2e == _T_153) begin
                                                                        mem_46 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h2f == wPos) begin
            mem_47 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h2f == _T_308) begin
                mem_47 <= _GEN_31;
              end else begin
                if (6'h2f == _T_303) begin
                  mem_47 <= _GEN_30;
                end else begin
                  if (6'h2f == _T_298) begin
                    mem_47 <= _GEN_29;
                  end else begin
                    if (6'h2f == _T_293) begin
                      mem_47 <= _GEN_28;
                    end else begin
                      if (6'h2f == _T_288) begin
                        mem_47 <= _GEN_27;
                      end else begin
                        if (6'h2f == _T_283) begin
                          mem_47 <= _GEN_26;
                        end else begin
                          if (6'h2f == _T_278) begin
                            mem_47 <= _GEN_25;
                          end else begin
                            if (6'h2f == _T_273) begin
                              mem_47 <= _GEN_24;
                            end else begin
                              if (6'h2f == _T_268) begin
                                mem_47 <= _GEN_23;
                              end else begin
                                if (6'h2f == _T_263) begin
                                  mem_47 <= _GEN_22;
                                end else begin
                                  if (6'h2f == _T_258) begin
                                    mem_47 <= _GEN_21;
                                  end else begin
                                    if (6'h2f == _T_253) begin
                                      mem_47 <= _GEN_20;
                                    end else begin
                                      if (6'h2f == _T_248) begin
                                        mem_47 <= _GEN_19;
                                      end else begin
                                        if (6'h2f == _T_243) begin
                                          mem_47 <= _GEN_18;
                                        end else begin
                                          if (6'h2f == _T_238) begin
                                            mem_47 <= _GEN_17;
                                          end else begin
                                            if (6'h2f == _T_233) begin
                                              mem_47 <= _GEN_16;
                                            end else begin
                                              if (6'h2f == _T_228) begin
                                                mem_47 <= _GEN_15;
                                              end else begin
                                                if (6'h2f == _T_223) begin
                                                  mem_47 <= _GEN_14;
                                                end else begin
                                                  if (6'h2f == _T_218) begin
                                                    mem_47 <= _GEN_13;
                                                  end else begin
                                                    if (6'h2f == _T_213) begin
                                                      mem_47 <= _GEN_12;
                                                    end else begin
                                                      if (6'h2f == _T_208) begin
                                                        mem_47 <= _GEN_11;
                                                      end else begin
                                                        if (6'h2f == _T_203) begin
                                                          mem_47 <= _GEN_10;
                                                        end else begin
                                                          if (6'h2f == _T_198) begin
                                                            mem_47 <= _GEN_9;
                                                          end else begin
                                                            if (6'h2f == _T_193) begin
                                                              mem_47 <= _GEN_8;
                                                            end else begin
                                                              if (6'h2f == _T_188) begin
                                                                mem_47 <= _GEN_7;
                                                              end else begin
                                                                if (6'h2f == _T_183) begin
                                                                  mem_47 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h2f == _T_178) begin
                                                                    mem_47 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h2f == _T_173) begin
                                                                      mem_47 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h2f == _T_168) begin
                                                                        mem_47 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h2f == _T_163) begin
                                                                          mem_47 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h2f == _T_158) begin
                                                                            mem_47 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h2f == _T_153) begin
                                                                              mem_47 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h2f == _T_308) begin
              mem_47 <= _GEN_31;
            end else begin
              if (6'h2f == _T_303) begin
                mem_47 <= _GEN_30;
              end else begin
                if (6'h2f == _T_298) begin
                  mem_47 <= _GEN_29;
                end else begin
                  if (6'h2f == _T_293) begin
                    mem_47 <= _GEN_28;
                  end else begin
                    if (6'h2f == _T_288) begin
                      mem_47 <= _GEN_27;
                    end else begin
                      if (6'h2f == _T_283) begin
                        mem_47 <= _GEN_26;
                      end else begin
                        if (6'h2f == _T_278) begin
                          mem_47 <= _GEN_25;
                        end else begin
                          if (6'h2f == _T_273) begin
                            mem_47 <= _GEN_24;
                          end else begin
                            if (6'h2f == _T_268) begin
                              mem_47 <= _GEN_23;
                            end else begin
                              if (6'h2f == _T_263) begin
                                mem_47 <= _GEN_22;
                              end else begin
                                if (6'h2f == _T_258) begin
                                  mem_47 <= _GEN_21;
                                end else begin
                                  if (6'h2f == _T_253) begin
                                    mem_47 <= _GEN_20;
                                  end else begin
                                    if (6'h2f == _T_248) begin
                                      mem_47 <= _GEN_19;
                                    end else begin
                                      if (6'h2f == _T_243) begin
                                        mem_47 <= _GEN_18;
                                      end else begin
                                        if (6'h2f == _T_238) begin
                                          mem_47 <= _GEN_17;
                                        end else begin
                                          if (6'h2f == _T_233) begin
                                            mem_47 <= _GEN_16;
                                          end else begin
                                            if (6'h2f == _T_228) begin
                                              mem_47 <= _GEN_15;
                                            end else begin
                                              if (6'h2f == _T_223) begin
                                                mem_47 <= _GEN_14;
                                              end else begin
                                                if (6'h2f == _T_218) begin
                                                  mem_47 <= _GEN_13;
                                                end else begin
                                                  if (6'h2f == _T_213) begin
                                                    mem_47 <= _GEN_12;
                                                  end else begin
                                                    if (6'h2f == _T_208) begin
                                                      mem_47 <= _GEN_11;
                                                    end else begin
                                                      if (6'h2f == _T_203) begin
                                                        mem_47 <= _GEN_10;
                                                      end else begin
                                                        if (6'h2f == _T_198) begin
                                                          mem_47 <= _GEN_9;
                                                        end else begin
                                                          if (6'h2f == _T_193) begin
                                                            mem_47 <= _GEN_8;
                                                          end else begin
                                                            if (6'h2f == _T_188) begin
                                                              mem_47 <= _GEN_7;
                                                            end else begin
                                                              if (6'h2f == _T_183) begin
                                                                mem_47 <= _GEN_6;
                                                              end else begin
                                                                if (6'h2f == _T_178) begin
                                                                  mem_47 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h2f == _T_173) begin
                                                                    mem_47 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h2f == _T_168) begin
                                                                      mem_47 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h2f == _T_163) begin
                                                                        mem_47 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h2f == _T_158) begin
                                                                          mem_47 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h2f == _T_153) begin
                                                                            mem_47 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h2f == _T_308) begin
            mem_47 <= _GEN_31;
          end else begin
            if (6'h2f == _T_303) begin
              mem_47 <= _GEN_30;
            end else begin
              if (6'h2f == _T_298) begin
                mem_47 <= _GEN_29;
              end else begin
                if (6'h2f == _T_293) begin
                  mem_47 <= _GEN_28;
                end else begin
                  if (6'h2f == _T_288) begin
                    mem_47 <= _GEN_27;
                  end else begin
                    if (6'h2f == _T_283) begin
                      mem_47 <= _GEN_26;
                    end else begin
                      if (6'h2f == _T_278) begin
                        mem_47 <= _GEN_25;
                      end else begin
                        if (6'h2f == _T_273) begin
                          mem_47 <= _GEN_24;
                        end else begin
                          if (6'h2f == _T_268) begin
                            mem_47 <= _GEN_23;
                          end else begin
                            if (6'h2f == _T_263) begin
                              mem_47 <= _GEN_22;
                            end else begin
                              if (6'h2f == _T_258) begin
                                mem_47 <= _GEN_21;
                              end else begin
                                if (6'h2f == _T_253) begin
                                  mem_47 <= _GEN_20;
                                end else begin
                                  if (6'h2f == _T_248) begin
                                    mem_47 <= _GEN_19;
                                  end else begin
                                    if (6'h2f == _T_243) begin
                                      mem_47 <= _GEN_18;
                                    end else begin
                                      if (6'h2f == _T_238) begin
                                        mem_47 <= _GEN_17;
                                      end else begin
                                        if (6'h2f == _T_233) begin
                                          mem_47 <= _GEN_16;
                                        end else begin
                                          if (6'h2f == _T_228) begin
                                            mem_47 <= _GEN_15;
                                          end else begin
                                            if (6'h2f == _T_223) begin
                                              mem_47 <= _GEN_14;
                                            end else begin
                                              if (6'h2f == _T_218) begin
                                                mem_47 <= _GEN_13;
                                              end else begin
                                                if (6'h2f == _T_213) begin
                                                  mem_47 <= _GEN_12;
                                                end else begin
                                                  if (6'h2f == _T_208) begin
                                                    mem_47 <= _GEN_11;
                                                  end else begin
                                                    if (6'h2f == _T_203) begin
                                                      mem_47 <= _GEN_10;
                                                    end else begin
                                                      if (6'h2f == _T_198) begin
                                                        mem_47 <= _GEN_9;
                                                      end else begin
                                                        if (6'h2f == _T_193) begin
                                                          mem_47 <= _GEN_8;
                                                        end else begin
                                                          if (6'h2f == _T_188) begin
                                                            mem_47 <= _GEN_7;
                                                          end else begin
                                                            if (6'h2f == _T_183) begin
                                                              mem_47 <= _GEN_6;
                                                            end else begin
                                                              if (6'h2f == _T_178) begin
                                                                mem_47 <= _GEN_5;
                                                              end else begin
                                                                if (6'h2f == _T_173) begin
                                                                  mem_47 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h2f == _T_168) begin
                                                                    mem_47 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h2f == _T_163) begin
                                                                      mem_47 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h2f == _T_158) begin
                                                                        mem_47 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h2f == _T_153) begin
                                                                          mem_47 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h2f == _T_308) begin
          mem_47 <= _GEN_31;
        end else begin
          if (6'h2f == _T_303) begin
            mem_47 <= _GEN_30;
          end else begin
            if (6'h2f == _T_298) begin
              mem_47 <= _GEN_29;
            end else begin
              if (6'h2f == _T_293) begin
                mem_47 <= _GEN_28;
              end else begin
                if (6'h2f == _T_288) begin
                  mem_47 <= _GEN_27;
                end else begin
                  if (6'h2f == _T_283) begin
                    mem_47 <= _GEN_26;
                  end else begin
                    if (6'h2f == _T_278) begin
                      mem_47 <= _GEN_25;
                    end else begin
                      if (6'h2f == _T_273) begin
                        mem_47 <= _GEN_24;
                      end else begin
                        if (6'h2f == _T_268) begin
                          mem_47 <= _GEN_23;
                        end else begin
                          if (6'h2f == _T_263) begin
                            mem_47 <= _GEN_22;
                          end else begin
                            if (6'h2f == _T_258) begin
                              mem_47 <= _GEN_21;
                            end else begin
                              if (6'h2f == _T_253) begin
                                mem_47 <= _GEN_20;
                              end else begin
                                if (6'h2f == _T_248) begin
                                  mem_47 <= _GEN_19;
                                end else begin
                                  if (6'h2f == _T_243) begin
                                    mem_47 <= _GEN_18;
                                  end else begin
                                    if (6'h2f == _T_238) begin
                                      mem_47 <= _GEN_17;
                                    end else begin
                                      if (6'h2f == _T_233) begin
                                        mem_47 <= _GEN_16;
                                      end else begin
                                        if (6'h2f == _T_228) begin
                                          mem_47 <= _GEN_15;
                                        end else begin
                                          if (6'h2f == _T_223) begin
                                            mem_47 <= _GEN_14;
                                          end else begin
                                            if (6'h2f == _T_218) begin
                                              mem_47 <= _GEN_13;
                                            end else begin
                                              if (6'h2f == _T_213) begin
                                                mem_47 <= _GEN_12;
                                              end else begin
                                                if (6'h2f == _T_208) begin
                                                  mem_47 <= _GEN_11;
                                                end else begin
                                                  if (6'h2f == _T_203) begin
                                                    mem_47 <= _GEN_10;
                                                  end else begin
                                                    if (6'h2f == _T_198) begin
                                                      mem_47 <= _GEN_9;
                                                    end else begin
                                                      if (6'h2f == _T_193) begin
                                                        mem_47 <= _GEN_8;
                                                      end else begin
                                                        if (6'h2f == _T_188) begin
                                                          mem_47 <= _GEN_7;
                                                        end else begin
                                                          if (6'h2f == _T_183) begin
                                                            mem_47 <= _GEN_6;
                                                          end else begin
                                                            if (6'h2f == _T_178) begin
                                                              mem_47 <= _GEN_5;
                                                            end else begin
                                                              if (6'h2f == _T_173) begin
                                                                mem_47 <= _GEN_4;
                                                              end else begin
                                                                if (6'h2f == _T_168) begin
                                                                  mem_47 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h2f == _T_163) begin
                                                                    mem_47 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h2f == _T_158) begin
                                                                      mem_47 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h2f == _T_153) begin
                                                                        mem_47 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h30 == wPos) begin
            mem_48 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h30 == _T_308) begin
                mem_48 <= _GEN_31;
              end else begin
                if (6'h30 == _T_303) begin
                  mem_48 <= _GEN_30;
                end else begin
                  if (6'h30 == _T_298) begin
                    mem_48 <= _GEN_29;
                  end else begin
                    if (6'h30 == _T_293) begin
                      mem_48 <= _GEN_28;
                    end else begin
                      if (6'h30 == _T_288) begin
                        mem_48 <= _GEN_27;
                      end else begin
                        if (6'h30 == _T_283) begin
                          mem_48 <= _GEN_26;
                        end else begin
                          if (6'h30 == _T_278) begin
                            mem_48 <= _GEN_25;
                          end else begin
                            if (6'h30 == _T_273) begin
                              mem_48 <= _GEN_24;
                            end else begin
                              if (6'h30 == _T_268) begin
                                mem_48 <= _GEN_23;
                              end else begin
                                if (6'h30 == _T_263) begin
                                  mem_48 <= _GEN_22;
                                end else begin
                                  if (6'h30 == _T_258) begin
                                    mem_48 <= _GEN_21;
                                  end else begin
                                    if (6'h30 == _T_253) begin
                                      mem_48 <= _GEN_20;
                                    end else begin
                                      if (6'h30 == _T_248) begin
                                        mem_48 <= _GEN_19;
                                      end else begin
                                        if (6'h30 == _T_243) begin
                                          mem_48 <= _GEN_18;
                                        end else begin
                                          if (6'h30 == _T_238) begin
                                            mem_48 <= _GEN_17;
                                          end else begin
                                            if (6'h30 == _T_233) begin
                                              mem_48 <= _GEN_16;
                                            end else begin
                                              if (6'h30 == _T_228) begin
                                                mem_48 <= _GEN_15;
                                              end else begin
                                                if (6'h30 == _T_223) begin
                                                  mem_48 <= _GEN_14;
                                                end else begin
                                                  if (6'h30 == _T_218) begin
                                                    mem_48 <= _GEN_13;
                                                  end else begin
                                                    if (6'h30 == _T_213) begin
                                                      mem_48 <= _GEN_12;
                                                    end else begin
                                                      if (6'h30 == _T_208) begin
                                                        mem_48 <= _GEN_11;
                                                      end else begin
                                                        if (6'h30 == _T_203) begin
                                                          mem_48 <= _GEN_10;
                                                        end else begin
                                                          if (6'h30 == _T_198) begin
                                                            mem_48 <= _GEN_9;
                                                          end else begin
                                                            if (6'h30 == _T_193) begin
                                                              mem_48 <= _GEN_8;
                                                            end else begin
                                                              if (6'h30 == _T_188) begin
                                                                mem_48 <= _GEN_7;
                                                              end else begin
                                                                if (6'h30 == _T_183) begin
                                                                  mem_48 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h30 == _T_178) begin
                                                                    mem_48 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h30 == _T_173) begin
                                                                      mem_48 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h30 == _T_168) begin
                                                                        mem_48 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h30 == _T_163) begin
                                                                          mem_48 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h30 == _T_158) begin
                                                                            mem_48 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h30 == _T_153) begin
                                                                              mem_48 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h30 == _T_308) begin
              mem_48 <= _GEN_31;
            end else begin
              if (6'h30 == _T_303) begin
                mem_48 <= _GEN_30;
              end else begin
                if (6'h30 == _T_298) begin
                  mem_48 <= _GEN_29;
                end else begin
                  if (6'h30 == _T_293) begin
                    mem_48 <= _GEN_28;
                  end else begin
                    if (6'h30 == _T_288) begin
                      mem_48 <= _GEN_27;
                    end else begin
                      if (6'h30 == _T_283) begin
                        mem_48 <= _GEN_26;
                      end else begin
                        if (6'h30 == _T_278) begin
                          mem_48 <= _GEN_25;
                        end else begin
                          if (6'h30 == _T_273) begin
                            mem_48 <= _GEN_24;
                          end else begin
                            if (6'h30 == _T_268) begin
                              mem_48 <= _GEN_23;
                            end else begin
                              if (6'h30 == _T_263) begin
                                mem_48 <= _GEN_22;
                              end else begin
                                if (6'h30 == _T_258) begin
                                  mem_48 <= _GEN_21;
                                end else begin
                                  if (6'h30 == _T_253) begin
                                    mem_48 <= _GEN_20;
                                  end else begin
                                    if (6'h30 == _T_248) begin
                                      mem_48 <= _GEN_19;
                                    end else begin
                                      if (6'h30 == _T_243) begin
                                        mem_48 <= _GEN_18;
                                      end else begin
                                        if (6'h30 == _T_238) begin
                                          mem_48 <= _GEN_17;
                                        end else begin
                                          if (6'h30 == _T_233) begin
                                            mem_48 <= _GEN_16;
                                          end else begin
                                            if (6'h30 == _T_228) begin
                                              mem_48 <= _GEN_15;
                                            end else begin
                                              if (6'h30 == _T_223) begin
                                                mem_48 <= _GEN_14;
                                              end else begin
                                                if (6'h30 == _T_218) begin
                                                  mem_48 <= _GEN_13;
                                                end else begin
                                                  if (6'h30 == _T_213) begin
                                                    mem_48 <= _GEN_12;
                                                  end else begin
                                                    if (6'h30 == _T_208) begin
                                                      mem_48 <= _GEN_11;
                                                    end else begin
                                                      if (6'h30 == _T_203) begin
                                                        mem_48 <= _GEN_10;
                                                      end else begin
                                                        if (6'h30 == _T_198) begin
                                                          mem_48 <= _GEN_9;
                                                        end else begin
                                                          if (6'h30 == _T_193) begin
                                                            mem_48 <= _GEN_8;
                                                          end else begin
                                                            if (6'h30 == _T_188) begin
                                                              mem_48 <= _GEN_7;
                                                            end else begin
                                                              if (6'h30 == _T_183) begin
                                                                mem_48 <= _GEN_6;
                                                              end else begin
                                                                if (6'h30 == _T_178) begin
                                                                  mem_48 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h30 == _T_173) begin
                                                                    mem_48 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h30 == _T_168) begin
                                                                      mem_48 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h30 == _T_163) begin
                                                                        mem_48 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h30 == _T_158) begin
                                                                          mem_48 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h30 == _T_153) begin
                                                                            mem_48 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h30 == _T_308) begin
            mem_48 <= _GEN_31;
          end else begin
            if (6'h30 == _T_303) begin
              mem_48 <= _GEN_30;
            end else begin
              if (6'h30 == _T_298) begin
                mem_48 <= _GEN_29;
              end else begin
                if (6'h30 == _T_293) begin
                  mem_48 <= _GEN_28;
                end else begin
                  if (6'h30 == _T_288) begin
                    mem_48 <= _GEN_27;
                  end else begin
                    if (6'h30 == _T_283) begin
                      mem_48 <= _GEN_26;
                    end else begin
                      if (6'h30 == _T_278) begin
                        mem_48 <= _GEN_25;
                      end else begin
                        if (6'h30 == _T_273) begin
                          mem_48 <= _GEN_24;
                        end else begin
                          if (6'h30 == _T_268) begin
                            mem_48 <= _GEN_23;
                          end else begin
                            if (6'h30 == _T_263) begin
                              mem_48 <= _GEN_22;
                            end else begin
                              if (6'h30 == _T_258) begin
                                mem_48 <= _GEN_21;
                              end else begin
                                if (6'h30 == _T_253) begin
                                  mem_48 <= _GEN_20;
                                end else begin
                                  if (6'h30 == _T_248) begin
                                    mem_48 <= _GEN_19;
                                  end else begin
                                    if (6'h30 == _T_243) begin
                                      mem_48 <= _GEN_18;
                                    end else begin
                                      if (6'h30 == _T_238) begin
                                        mem_48 <= _GEN_17;
                                      end else begin
                                        if (6'h30 == _T_233) begin
                                          mem_48 <= _GEN_16;
                                        end else begin
                                          if (6'h30 == _T_228) begin
                                            mem_48 <= _GEN_15;
                                          end else begin
                                            if (6'h30 == _T_223) begin
                                              mem_48 <= _GEN_14;
                                            end else begin
                                              if (6'h30 == _T_218) begin
                                                mem_48 <= _GEN_13;
                                              end else begin
                                                if (6'h30 == _T_213) begin
                                                  mem_48 <= _GEN_12;
                                                end else begin
                                                  if (6'h30 == _T_208) begin
                                                    mem_48 <= _GEN_11;
                                                  end else begin
                                                    if (6'h30 == _T_203) begin
                                                      mem_48 <= _GEN_10;
                                                    end else begin
                                                      if (6'h30 == _T_198) begin
                                                        mem_48 <= _GEN_9;
                                                      end else begin
                                                        if (6'h30 == _T_193) begin
                                                          mem_48 <= _GEN_8;
                                                        end else begin
                                                          if (6'h30 == _T_188) begin
                                                            mem_48 <= _GEN_7;
                                                          end else begin
                                                            if (6'h30 == _T_183) begin
                                                              mem_48 <= _GEN_6;
                                                            end else begin
                                                              if (6'h30 == _T_178) begin
                                                                mem_48 <= _GEN_5;
                                                              end else begin
                                                                if (6'h30 == _T_173) begin
                                                                  mem_48 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h30 == _T_168) begin
                                                                    mem_48 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h30 == _T_163) begin
                                                                      mem_48 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h30 == _T_158) begin
                                                                        mem_48 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h30 == _T_153) begin
                                                                          mem_48 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h30 == _T_308) begin
          mem_48 <= _GEN_31;
        end else begin
          if (6'h30 == _T_303) begin
            mem_48 <= _GEN_30;
          end else begin
            if (6'h30 == _T_298) begin
              mem_48 <= _GEN_29;
            end else begin
              if (6'h30 == _T_293) begin
                mem_48 <= _GEN_28;
              end else begin
                if (6'h30 == _T_288) begin
                  mem_48 <= _GEN_27;
                end else begin
                  if (6'h30 == _T_283) begin
                    mem_48 <= _GEN_26;
                  end else begin
                    if (6'h30 == _T_278) begin
                      mem_48 <= _GEN_25;
                    end else begin
                      if (6'h30 == _T_273) begin
                        mem_48 <= _GEN_24;
                      end else begin
                        if (6'h30 == _T_268) begin
                          mem_48 <= _GEN_23;
                        end else begin
                          if (6'h30 == _T_263) begin
                            mem_48 <= _GEN_22;
                          end else begin
                            if (6'h30 == _T_258) begin
                              mem_48 <= _GEN_21;
                            end else begin
                              if (6'h30 == _T_253) begin
                                mem_48 <= _GEN_20;
                              end else begin
                                if (6'h30 == _T_248) begin
                                  mem_48 <= _GEN_19;
                                end else begin
                                  if (6'h30 == _T_243) begin
                                    mem_48 <= _GEN_18;
                                  end else begin
                                    if (6'h30 == _T_238) begin
                                      mem_48 <= _GEN_17;
                                    end else begin
                                      if (6'h30 == _T_233) begin
                                        mem_48 <= _GEN_16;
                                      end else begin
                                        if (6'h30 == _T_228) begin
                                          mem_48 <= _GEN_15;
                                        end else begin
                                          if (6'h30 == _T_223) begin
                                            mem_48 <= _GEN_14;
                                          end else begin
                                            if (6'h30 == _T_218) begin
                                              mem_48 <= _GEN_13;
                                            end else begin
                                              if (6'h30 == _T_213) begin
                                                mem_48 <= _GEN_12;
                                              end else begin
                                                if (6'h30 == _T_208) begin
                                                  mem_48 <= _GEN_11;
                                                end else begin
                                                  if (6'h30 == _T_203) begin
                                                    mem_48 <= _GEN_10;
                                                  end else begin
                                                    if (6'h30 == _T_198) begin
                                                      mem_48 <= _GEN_9;
                                                    end else begin
                                                      if (6'h30 == _T_193) begin
                                                        mem_48 <= _GEN_8;
                                                      end else begin
                                                        if (6'h30 == _T_188) begin
                                                          mem_48 <= _GEN_7;
                                                        end else begin
                                                          if (6'h30 == _T_183) begin
                                                            mem_48 <= _GEN_6;
                                                          end else begin
                                                            if (6'h30 == _T_178) begin
                                                              mem_48 <= _GEN_5;
                                                            end else begin
                                                              if (6'h30 == _T_173) begin
                                                                mem_48 <= _GEN_4;
                                                              end else begin
                                                                if (6'h30 == _T_168) begin
                                                                  mem_48 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h30 == _T_163) begin
                                                                    mem_48 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h30 == _T_158) begin
                                                                      mem_48 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h30 == _T_153) begin
                                                                        mem_48 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h31 == wPos) begin
            mem_49 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h31 == _T_308) begin
                mem_49 <= _GEN_31;
              end else begin
                if (6'h31 == _T_303) begin
                  mem_49 <= _GEN_30;
                end else begin
                  if (6'h31 == _T_298) begin
                    mem_49 <= _GEN_29;
                  end else begin
                    if (6'h31 == _T_293) begin
                      mem_49 <= _GEN_28;
                    end else begin
                      if (6'h31 == _T_288) begin
                        mem_49 <= _GEN_27;
                      end else begin
                        if (6'h31 == _T_283) begin
                          mem_49 <= _GEN_26;
                        end else begin
                          if (6'h31 == _T_278) begin
                            mem_49 <= _GEN_25;
                          end else begin
                            if (6'h31 == _T_273) begin
                              mem_49 <= _GEN_24;
                            end else begin
                              if (6'h31 == _T_268) begin
                                mem_49 <= _GEN_23;
                              end else begin
                                if (6'h31 == _T_263) begin
                                  mem_49 <= _GEN_22;
                                end else begin
                                  if (6'h31 == _T_258) begin
                                    mem_49 <= _GEN_21;
                                  end else begin
                                    if (6'h31 == _T_253) begin
                                      mem_49 <= _GEN_20;
                                    end else begin
                                      if (6'h31 == _T_248) begin
                                        mem_49 <= _GEN_19;
                                      end else begin
                                        if (6'h31 == _T_243) begin
                                          mem_49 <= _GEN_18;
                                        end else begin
                                          if (6'h31 == _T_238) begin
                                            mem_49 <= _GEN_17;
                                          end else begin
                                            if (6'h31 == _T_233) begin
                                              mem_49 <= _GEN_16;
                                            end else begin
                                              if (6'h31 == _T_228) begin
                                                mem_49 <= _GEN_15;
                                              end else begin
                                                if (6'h31 == _T_223) begin
                                                  mem_49 <= _GEN_14;
                                                end else begin
                                                  if (6'h31 == _T_218) begin
                                                    mem_49 <= _GEN_13;
                                                  end else begin
                                                    if (6'h31 == _T_213) begin
                                                      mem_49 <= _GEN_12;
                                                    end else begin
                                                      if (6'h31 == _T_208) begin
                                                        mem_49 <= _GEN_11;
                                                      end else begin
                                                        if (6'h31 == _T_203) begin
                                                          mem_49 <= _GEN_10;
                                                        end else begin
                                                          if (6'h31 == _T_198) begin
                                                            mem_49 <= _GEN_9;
                                                          end else begin
                                                            if (6'h31 == _T_193) begin
                                                              mem_49 <= _GEN_8;
                                                            end else begin
                                                              if (6'h31 == _T_188) begin
                                                                mem_49 <= _GEN_7;
                                                              end else begin
                                                                if (6'h31 == _T_183) begin
                                                                  mem_49 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h31 == _T_178) begin
                                                                    mem_49 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h31 == _T_173) begin
                                                                      mem_49 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h31 == _T_168) begin
                                                                        mem_49 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h31 == _T_163) begin
                                                                          mem_49 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h31 == _T_158) begin
                                                                            mem_49 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h31 == _T_153) begin
                                                                              mem_49 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h31 == _T_308) begin
              mem_49 <= _GEN_31;
            end else begin
              if (6'h31 == _T_303) begin
                mem_49 <= _GEN_30;
              end else begin
                if (6'h31 == _T_298) begin
                  mem_49 <= _GEN_29;
                end else begin
                  if (6'h31 == _T_293) begin
                    mem_49 <= _GEN_28;
                  end else begin
                    if (6'h31 == _T_288) begin
                      mem_49 <= _GEN_27;
                    end else begin
                      if (6'h31 == _T_283) begin
                        mem_49 <= _GEN_26;
                      end else begin
                        if (6'h31 == _T_278) begin
                          mem_49 <= _GEN_25;
                        end else begin
                          if (6'h31 == _T_273) begin
                            mem_49 <= _GEN_24;
                          end else begin
                            if (6'h31 == _T_268) begin
                              mem_49 <= _GEN_23;
                            end else begin
                              if (6'h31 == _T_263) begin
                                mem_49 <= _GEN_22;
                              end else begin
                                if (6'h31 == _T_258) begin
                                  mem_49 <= _GEN_21;
                                end else begin
                                  if (6'h31 == _T_253) begin
                                    mem_49 <= _GEN_20;
                                  end else begin
                                    if (6'h31 == _T_248) begin
                                      mem_49 <= _GEN_19;
                                    end else begin
                                      if (6'h31 == _T_243) begin
                                        mem_49 <= _GEN_18;
                                      end else begin
                                        if (6'h31 == _T_238) begin
                                          mem_49 <= _GEN_17;
                                        end else begin
                                          if (6'h31 == _T_233) begin
                                            mem_49 <= _GEN_16;
                                          end else begin
                                            if (6'h31 == _T_228) begin
                                              mem_49 <= _GEN_15;
                                            end else begin
                                              if (6'h31 == _T_223) begin
                                                mem_49 <= _GEN_14;
                                              end else begin
                                                if (6'h31 == _T_218) begin
                                                  mem_49 <= _GEN_13;
                                                end else begin
                                                  if (6'h31 == _T_213) begin
                                                    mem_49 <= _GEN_12;
                                                  end else begin
                                                    if (6'h31 == _T_208) begin
                                                      mem_49 <= _GEN_11;
                                                    end else begin
                                                      if (6'h31 == _T_203) begin
                                                        mem_49 <= _GEN_10;
                                                      end else begin
                                                        if (6'h31 == _T_198) begin
                                                          mem_49 <= _GEN_9;
                                                        end else begin
                                                          if (6'h31 == _T_193) begin
                                                            mem_49 <= _GEN_8;
                                                          end else begin
                                                            if (6'h31 == _T_188) begin
                                                              mem_49 <= _GEN_7;
                                                            end else begin
                                                              if (6'h31 == _T_183) begin
                                                                mem_49 <= _GEN_6;
                                                              end else begin
                                                                if (6'h31 == _T_178) begin
                                                                  mem_49 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h31 == _T_173) begin
                                                                    mem_49 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h31 == _T_168) begin
                                                                      mem_49 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h31 == _T_163) begin
                                                                        mem_49 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h31 == _T_158) begin
                                                                          mem_49 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h31 == _T_153) begin
                                                                            mem_49 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h31 == _T_308) begin
            mem_49 <= _GEN_31;
          end else begin
            if (6'h31 == _T_303) begin
              mem_49 <= _GEN_30;
            end else begin
              if (6'h31 == _T_298) begin
                mem_49 <= _GEN_29;
              end else begin
                if (6'h31 == _T_293) begin
                  mem_49 <= _GEN_28;
                end else begin
                  if (6'h31 == _T_288) begin
                    mem_49 <= _GEN_27;
                  end else begin
                    if (6'h31 == _T_283) begin
                      mem_49 <= _GEN_26;
                    end else begin
                      if (6'h31 == _T_278) begin
                        mem_49 <= _GEN_25;
                      end else begin
                        if (6'h31 == _T_273) begin
                          mem_49 <= _GEN_24;
                        end else begin
                          if (6'h31 == _T_268) begin
                            mem_49 <= _GEN_23;
                          end else begin
                            if (6'h31 == _T_263) begin
                              mem_49 <= _GEN_22;
                            end else begin
                              if (6'h31 == _T_258) begin
                                mem_49 <= _GEN_21;
                              end else begin
                                if (6'h31 == _T_253) begin
                                  mem_49 <= _GEN_20;
                                end else begin
                                  if (6'h31 == _T_248) begin
                                    mem_49 <= _GEN_19;
                                  end else begin
                                    if (6'h31 == _T_243) begin
                                      mem_49 <= _GEN_18;
                                    end else begin
                                      if (6'h31 == _T_238) begin
                                        mem_49 <= _GEN_17;
                                      end else begin
                                        if (6'h31 == _T_233) begin
                                          mem_49 <= _GEN_16;
                                        end else begin
                                          if (6'h31 == _T_228) begin
                                            mem_49 <= _GEN_15;
                                          end else begin
                                            if (6'h31 == _T_223) begin
                                              mem_49 <= _GEN_14;
                                            end else begin
                                              if (6'h31 == _T_218) begin
                                                mem_49 <= _GEN_13;
                                              end else begin
                                                if (6'h31 == _T_213) begin
                                                  mem_49 <= _GEN_12;
                                                end else begin
                                                  if (6'h31 == _T_208) begin
                                                    mem_49 <= _GEN_11;
                                                  end else begin
                                                    if (6'h31 == _T_203) begin
                                                      mem_49 <= _GEN_10;
                                                    end else begin
                                                      if (6'h31 == _T_198) begin
                                                        mem_49 <= _GEN_9;
                                                      end else begin
                                                        if (6'h31 == _T_193) begin
                                                          mem_49 <= _GEN_8;
                                                        end else begin
                                                          if (6'h31 == _T_188) begin
                                                            mem_49 <= _GEN_7;
                                                          end else begin
                                                            if (6'h31 == _T_183) begin
                                                              mem_49 <= _GEN_6;
                                                            end else begin
                                                              if (6'h31 == _T_178) begin
                                                                mem_49 <= _GEN_5;
                                                              end else begin
                                                                if (6'h31 == _T_173) begin
                                                                  mem_49 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h31 == _T_168) begin
                                                                    mem_49 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h31 == _T_163) begin
                                                                      mem_49 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h31 == _T_158) begin
                                                                        mem_49 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h31 == _T_153) begin
                                                                          mem_49 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h31 == _T_308) begin
          mem_49 <= _GEN_31;
        end else begin
          if (6'h31 == _T_303) begin
            mem_49 <= _GEN_30;
          end else begin
            if (6'h31 == _T_298) begin
              mem_49 <= _GEN_29;
            end else begin
              if (6'h31 == _T_293) begin
                mem_49 <= _GEN_28;
              end else begin
                if (6'h31 == _T_288) begin
                  mem_49 <= _GEN_27;
                end else begin
                  if (6'h31 == _T_283) begin
                    mem_49 <= _GEN_26;
                  end else begin
                    if (6'h31 == _T_278) begin
                      mem_49 <= _GEN_25;
                    end else begin
                      if (6'h31 == _T_273) begin
                        mem_49 <= _GEN_24;
                      end else begin
                        if (6'h31 == _T_268) begin
                          mem_49 <= _GEN_23;
                        end else begin
                          if (6'h31 == _T_263) begin
                            mem_49 <= _GEN_22;
                          end else begin
                            if (6'h31 == _T_258) begin
                              mem_49 <= _GEN_21;
                            end else begin
                              if (6'h31 == _T_253) begin
                                mem_49 <= _GEN_20;
                              end else begin
                                if (6'h31 == _T_248) begin
                                  mem_49 <= _GEN_19;
                                end else begin
                                  if (6'h31 == _T_243) begin
                                    mem_49 <= _GEN_18;
                                  end else begin
                                    if (6'h31 == _T_238) begin
                                      mem_49 <= _GEN_17;
                                    end else begin
                                      if (6'h31 == _T_233) begin
                                        mem_49 <= _GEN_16;
                                      end else begin
                                        if (6'h31 == _T_228) begin
                                          mem_49 <= _GEN_15;
                                        end else begin
                                          if (6'h31 == _T_223) begin
                                            mem_49 <= _GEN_14;
                                          end else begin
                                            if (6'h31 == _T_218) begin
                                              mem_49 <= _GEN_13;
                                            end else begin
                                              if (6'h31 == _T_213) begin
                                                mem_49 <= _GEN_12;
                                              end else begin
                                                if (6'h31 == _T_208) begin
                                                  mem_49 <= _GEN_11;
                                                end else begin
                                                  if (6'h31 == _T_203) begin
                                                    mem_49 <= _GEN_10;
                                                  end else begin
                                                    if (6'h31 == _T_198) begin
                                                      mem_49 <= _GEN_9;
                                                    end else begin
                                                      if (6'h31 == _T_193) begin
                                                        mem_49 <= _GEN_8;
                                                      end else begin
                                                        if (6'h31 == _T_188) begin
                                                          mem_49 <= _GEN_7;
                                                        end else begin
                                                          if (6'h31 == _T_183) begin
                                                            mem_49 <= _GEN_6;
                                                          end else begin
                                                            if (6'h31 == _T_178) begin
                                                              mem_49 <= _GEN_5;
                                                            end else begin
                                                              if (6'h31 == _T_173) begin
                                                                mem_49 <= _GEN_4;
                                                              end else begin
                                                                if (6'h31 == _T_168) begin
                                                                  mem_49 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h31 == _T_163) begin
                                                                    mem_49 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h31 == _T_158) begin
                                                                      mem_49 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h31 == _T_153) begin
                                                                        mem_49 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h32 == wPos) begin
            mem_50 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h32 == _T_308) begin
                mem_50 <= _GEN_31;
              end else begin
                if (6'h32 == _T_303) begin
                  mem_50 <= _GEN_30;
                end else begin
                  if (6'h32 == _T_298) begin
                    mem_50 <= _GEN_29;
                  end else begin
                    if (6'h32 == _T_293) begin
                      mem_50 <= _GEN_28;
                    end else begin
                      if (6'h32 == _T_288) begin
                        mem_50 <= _GEN_27;
                      end else begin
                        if (6'h32 == _T_283) begin
                          mem_50 <= _GEN_26;
                        end else begin
                          if (6'h32 == _T_278) begin
                            mem_50 <= _GEN_25;
                          end else begin
                            if (6'h32 == _T_273) begin
                              mem_50 <= _GEN_24;
                            end else begin
                              if (6'h32 == _T_268) begin
                                mem_50 <= _GEN_23;
                              end else begin
                                if (6'h32 == _T_263) begin
                                  mem_50 <= _GEN_22;
                                end else begin
                                  if (6'h32 == _T_258) begin
                                    mem_50 <= _GEN_21;
                                  end else begin
                                    if (6'h32 == _T_253) begin
                                      mem_50 <= _GEN_20;
                                    end else begin
                                      if (6'h32 == _T_248) begin
                                        mem_50 <= _GEN_19;
                                      end else begin
                                        if (6'h32 == _T_243) begin
                                          mem_50 <= _GEN_18;
                                        end else begin
                                          if (6'h32 == _T_238) begin
                                            mem_50 <= _GEN_17;
                                          end else begin
                                            if (6'h32 == _T_233) begin
                                              mem_50 <= _GEN_16;
                                            end else begin
                                              if (6'h32 == _T_228) begin
                                                mem_50 <= _GEN_15;
                                              end else begin
                                                if (6'h32 == _T_223) begin
                                                  mem_50 <= _GEN_14;
                                                end else begin
                                                  if (6'h32 == _T_218) begin
                                                    mem_50 <= _GEN_13;
                                                  end else begin
                                                    if (6'h32 == _T_213) begin
                                                      mem_50 <= _GEN_12;
                                                    end else begin
                                                      if (6'h32 == _T_208) begin
                                                        mem_50 <= _GEN_11;
                                                      end else begin
                                                        if (6'h32 == _T_203) begin
                                                          mem_50 <= _GEN_10;
                                                        end else begin
                                                          if (6'h32 == _T_198) begin
                                                            mem_50 <= _GEN_9;
                                                          end else begin
                                                            if (6'h32 == _T_193) begin
                                                              mem_50 <= _GEN_8;
                                                            end else begin
                                                              if (6'h32 == _T_188) begin
                                                                mem_50 <= _GEN_7;
                                                              end else begin
                                                                if (6'h32 == _T_183) begin
                                                                  mem_50 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h32 == _T_178) begin
                                                                    mem_50 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h32 == _T_173) begin
                                                                      mem_50 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h32 == _T_168) begin
                                                                        mem_50 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h32 == _T_163) begin
                                                                          mem_50 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h32 == _T_158) begin
                                                                            mem_50 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h32 == _T_153) begin
                                                                              mem_50 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h32 == _T_308) begin
              mem_50 <= _GEN_31;
            end else begin
              if (6'h32 == _T_303) begin
                mem_50 <= _GEN_30;
              end else begin
                if (6'h32 == _T_298) begin
                  mem_50 <= _GEN_29;
                end else begin
                  if (6'h32 == _T_293) begin
                    mem_50 <= _GEN_28;
                  end else begin
                    if (6'h32 == _T_288) begin
                      mem_50 <= _GEN_27;
                    end else begin
                      if (6'h32 == _T_283) begin
                        mem_50 <= _GEN_26;
                      end else begin
                        if (6'h32 == _T_278) begin
                          mem_50 <= _GEN_25;
                        end else begin
                          if (6'h32 == _T_273) begin
                            mem_50 <= _GEN_24;
                          end else begin
                            if (6'h32 == _T_268) begin
                              mem_50 <= _GEN_23;
                            end else begin
                              if (6'h32 == _T_263) begin
                                mem_50 <= _GEN_22;
                              end else begin
                                if (6'h32 == _T_258) begin
                                  mem_50 <= _GEN_21;
                                end else begin
                                  if (6'h32 == _T_253) begin
                                    mem_50 <= _GEN_20;
                                  end else begin
                                    if (6'h32 == _T_248) begin
                                      mem_50 <= _GEN_19;
                                    end else begin
                                      if (6'h32 == _T_243) begin
                                        mem_50 <= _GEN_18;
                                      end else begin
                                        if (6'h32 == _T_238) begin
                                          mem_50 <= _GEN_17;
                                        end else begin
                                          if (6'h32 == _T_233) begin
                                            mem_50 <= _GEN_16;
                                          end else begin
                                            if (6'h32 == _T_228) begin
                                              mem_50 <= _GEN_15;
                                            end else begin
                                              if (6'h32 == _T_223) begin
                                                mem_50 <= _GEN_14;
                                              end else begin
                                                if (6'h32 == _T_218) begin
                                                  mem_50 <= _GEN_13;
                                                end else begin
                                                  if (6'h32 == _T_213) begin
                                                    mem_50 <= _GEN_12;
                                                  end else begin
                                                    if (6'h32 == _T_208) begin
                                                      mem_50 <= _GEN_11;
                                                    end else begin
                                                      if (6'h32 == _T_203) begin
                                                        mem_50 <= _GEN_10;
                                                      end else begin
                                                        if (6'h32 == _T_198) begin
                                                          mem_50 <= _GEN_9;
                                                        end else begin
                                                          if (6'h32 == _T_193) begin
                                                            mem_50 <= _GEN_8;
                                                          end else begin
                                                            if (6'h32 == _T_188) begin
                                                              mem_50 <= _GEN_7;
                                                            end else begin
                                                              if (6'h32 == _T_183) begin
                                                                mem_50 <= _GEN_6;
                                                              end else begin
                                                                if (6'h32 == _T_178) begin
                                                                  mem_50 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h32 == _T_173) begin
                                                                    mem_50 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h32 == _T_168) begin
                                                                      mem_50 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h32 == _T_163) begin
                                                                        mem_50 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h32 == _T_158) begin
                                                                          mem_50 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h32 == _T_153) begin
                                                                            mem_50 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h32 == _T_308) begin
            mem_50 <= _GEN_31;
          end else begin
            if (6'h32 == _T_303) begin
              mem_50 <= _GEN_30;
            end else begin
              if (6'h32 == _T_298) begin
                mem_50 <= _GEN_29;
              end else begin
                if (6'h32 == _T_293) begin
                  mem_50 <= _GEN_28;
                end else begin
                  if (6'h32 == _T_288) begin
                    mem_50 <= _GEN_27;
                  end else begin
                    if (6'h32 == _T_283) begin
                      mem_50 <= _GEN_26;
                    end else begin
                      if (6'h32 == _T_278) begin
                        mem_50 <= _GEN_25;
                      end else begin
                        if (6'h32 == _T_273) begin
                          mem_50 <= _GEN_24;
                        end else begin
                          if (6'h32 == _T_268) begin
                            mem_50 <= _GEN_23;
                          end else begin
                            if (6'h32 == _T_263) begin
                              mem_50 <= _GEN_22;
                            end else begin
                              if (6'h32 == _T_258) begin
                                mem_50 <= _GEN_21;
                              end else begin
                                if (6'h32 == _T_253) begin
                                  mem_50 <= _GEN_20;
                                end else begin
                                  if (6'h32 == _T_248) begin
                                    mem_50 <= _GEN_19;
                                  end else begin
                                    if (6'h32 == _T_243) begin
                                      mem_50 <= _GEN_18;
                                    end else begin
                                      if (6'h32 == _T_238) begin
                                        mem_50 <= _GEN_17;
                                      end else begin
                                        if (6'h32 == _T_233) begin
                                          mem_50 <= _GEN_16;
                                        end else begin
                                          if (6'h32 == _T_228) begin
                                            mem_50 <= _GEN_15;
                                          end else begin
                                            if (6'h32 == _T_223) begin
                                              mem_50 <= _GEN_14;
                                            end else begin
                                              if (6'h32 == _T_218) begin
                                                mem_50 <= _GEN_13;
                                              end else begin
                                                if (6'h32 == _T_213) begin
                                                  mem_50 <= _GEN_12;
                                                end else begin
                                                  if (6'h32 == _T_208) begin
                                                    mem_50 <= _GEN_11;
                                                  end else begin
                                                    if (6'h32 == _T_203) begin
                                                      mem_50 <= _GEN_10;
                                                    end else begin
                                                      if (6'h32 == _T_198) begin
                                                        mem_50 <= _GEN_9;
                                                      end else begin
                                                        if (6'h32 == _T_193) begin
                                                          mem_50 <= _GEN_8;
                                                        end else begin
                                                          if (6'h32 == _T_188) begin
                                                            mem_50 <= _GEN_7;
                                                          end else begin
                                                            if (6'h32 == _T_183) begin
                                                              mem_50 <= _GEN_6;
                                                            end else begin
                                                              if (6'h32 == _T_178) begin
                                                                mem_50 <= _GEN_5;
                                                              end else begin
                                                                if (6'h32 == _T_173) begin
                                                                  mem_50 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h32 == _T_168) begin
                                                                    mem_50 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h32 == _T_163) begin
                                                                      mem_50 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h32 == _T_158) begin
                                                                        mem_50 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h32 == _T_153) begin
                                                                          mem_50 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h32 == _T_308) begin
          mem_50 <= _GEN_31;
        end else begin
          if (6'h32 == _T_303) begin
            mem_50 <= _GEN_30;
          end else begin
            if (6'h32 == _T_298) begin
              mem_50 <= _GEN_29;
            end else begin
              if (6'h32 == _T_293) begin
                mem_50 <= _GEN_28;
              end else begin
                if (6'h32 == _T_288) begin
                  mem_50 <= _GEN_27;
                end else begin
                  if (6'h32 == _T_283) begin
                    mem_50 <= _GEN_26;
                  end else begin
                    if (6'h32 == _T_278) begin
                      mem_50 <= _GEN_25;
                    end else begin
                      if (6'h32 == _T_273) begin
                        mem_50 <= _GEN_24;
                      end else begin
                        if (6'h32 == _T_268) begin
                          mem_50 <= _GEN_23;
                        end else begin
                          if (6'h32 == _T_263) begin
                            mem_50 <= _GEN_22;
                          end else begin
                            if (6'h32 == _T_258) begin
                              mem_50 <= _GEN_21;
                            end else begin
                              if (6'h32 == _T_253) begin
                                mem_50 <= _GEN_20;
                              end else begin
                                if (6'h32 == _T_248) begin
                                  mem_50 <= _GEN_19;
                                end else begin
                                  if (6'h32 == _T_243) begin
                                    mem_50 <= _GEN_18;
                                  end else begin
                                    if (6'h32 == _T_238) begin
                                      mem_50 <= _GEN_17;
                                    end else begin
                                      if (6'h32 == _T_233) begin
                                        mem_50 <= _GEN_16;
                                      end else begin
                                        if (6'h32 == _T_228) begin
                                          mem_50 <= _GEN_15;
                                        end else begin
                                          if (6'h32 == _T_223) begin
                                            mem_50 <= _GEN_14;
                                          end else begin
                                            if (6'h32 == _T_218) begin
                                              mem_50 <= _GEN_13;
                                            end else begin
                                              if (6'h32 == _T_213) begin
                                                mem_50 <= _GEN_12;
                                              end else begin
                                                if (6'h32 == _T_208) begin
                                                  mem_50 <= _GEN_11;
                                                end else begin
                                                  if (6'h32 == _T_203) begin
                                                    mem_50 <= _GEN_10;
                                                  end else begin
                                                    if (6'h32 == _T_198) begin
                                                      mem_50 <= _GEN_9;
                                                    end else begin
                                                      if (6'h32 == _T_193) begin
                                                        mem_50 <= _GEN_8;
                                                      end else begin
                                                        if (6'h32 == _T_188) begin
                                                          mem_50 <= _GEN_7;
                                                        end else begin
                                                          if (6'h32 == _T_183) begin
                                                            mem_50 <= _GEN_6;
                                                          end else begin
                                                            if (6'h32 == _T_178) begin
                                                              mem_50 <= _GEN_5;
                                                            end else begin
                                                              if (6'h32 == _T_173) begin
                                                                mem_50 <= _GEN_4;
                                                              end else begin
                                                                if (6'h32 == _T_168) begin
                                                                  mem_50 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h32 == _T_163) begin
                                                                    mem_50 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h32 == _T_158) begin
                                                                      mem_50 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h32 == _T_153) begin
                                                                        mem_50 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h33 == wPos) begin
            mem_51 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h33 == _T_308) begin
                mem_51 <= _GEN_31;
              end else begin
                if (6'h33 == _T_303) begin
                  mem_51 <= _GEN_30;
                end else begin
                  if (6'h33 == _T_298) begin
                    mem_51 <= _GEN_29;
                  end else begin
                    if (6'h33 == _T_293) begin
                      mem_51 <= _GEN_28;
                    end else begin
                      if (6'h33 == _T_288) begin
                        mem_51 <= _GEN_27;
                      end else begin
                        if (6'h33 == _T_283) begin
                          mem_51 <= _GEN_26;
                        end else begin
                          if (6'h33 == _T_278) begin
                            mem_51 <= _GEN_25;
                          end else begin
                            if (6'h33 == _T_273) begin
                              mem_51 <= _GEN_24;
                            end else begin
                              if (6'h33 == _T_268) begin
                                mem_51 <= _GEN_23;
                              end else begin
                                if (6'h33 == _T_263) begin
                                  mem_51 <= _GEN_22;
                                end else begin
                                  if (6'h33 == _T_258) begin
                                    mem_51 <= _GEN_21;
                                  end else begin
                                    if (6'h33 == _T_253) begin
                                      mem_51 <= _GEN_20;
                                    end else begin
                                      if (6'h33 == _T_248) begin
                                        mem_51 <= _GEN_19;
                                      end else begin
                                        if (6'h33 == _T_243) begin
                                          mem_51 <= _GEN_18;
                                        end else begin
                                          if (6'h33 == _T_238) begin
                                            mem_51 <= _GEN_17;
                                          end else begin
                                            if (6'h33 == _T_233) begin
                                              mem_51 <= _GEN_16;
                                            end else begin
                                              if (6'h33 == _T_228) begin
                                                mem_51 <= _GEN_15;
                                              end else begin
                                                if (6'h33 == _T_223) begin
                                                  mem_51 <= _GEN_14;
                                                end else begin
                                                  if (6'h33 == _T_218) begin
                                                    mem_51 <= _GEN_13;
                                                  end else begin
                                                    if (6'h33 == _T_213) begin
                                                      mem_51 <= _GEN_12;
                                                    end else begin
                                                      if (6'h33 == _T_208) begin
                                                        mem_51 <= _GEN_11;
                                                      end else begin
                                                        if (6'h33 == _T_203) begin
                                                          mem_51 <= _GEN_10;
                                                        end else begin
                                                          if (6'h33 == _T_198) begin
                                                            mem_51 <= _GEN_9;
                                                          end else begin
                                                            if (6'h33 == _T_193) begin
                                                              mem_51 <= _GEN_8;
                                                            end else begin
                                                              if (6'h33 == _T_188) begin
                                                                mem_51 <= _GEN_7;
                                                              end else begin
                                                                if (6'h33 == _T_183) begin
                                                                  mem_51 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h33 == _T_178) begin
                                                                    mem_51 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h33 == _T_173) begin
                                                                      mem_51 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h33 == _T_168) begin
                                                                        mem_51 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h33 == _T_163) begin
                                                                          mem_51 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h33 == _T_158) begin
                                                                            mem_51 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h33 == _T_153) begin
                                                                              mem_51 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h33 == _T_308) begin
              mem_51 <= _GEN_31;
            end else begin
              if (6'h33 == _T_303) begin
                mem_51 <= _GEN_30;
              end else begin
                if (6'h33 == _T_298) begin
                  mem_51 <= _GEN_29;
                end else begin
                  if (6'h33 == _T_293) begin
                    mem_51 <= _GEN_28;
                  end else begin
                    if (6'h33 == _T_288) begin
                      mem_51 <= _GEN_27;
                    end else begin
                      if (6'h33 == _T_283) begin
                        mem_51 <= _GEN_26;
                      end else begin
                        if (6'h33 == _T_278) begin
                          mem_51 <= _GEN_25;
                        end else begin
                          if (6'h33 == _T_273) begin
                            mem_51 <= _GEN_24;
                          end else begin
                            if (6'h33 == _T_268) begin
                              mem_51 <= _GEN_23;
                            end else begin
                              if (6'h33 == _T_263) begin
                                mem_51 <= _GEN_22;
                              end else begin
                                if (6'h33 == _T_258) begin
                                  mem_51 <= _GEN_21;
                                end else begin
                                  if (6'h33 == _T_253) begin
                                    mem_51 <= _GEN_20;
                                  end else begin
                                    if (6'h33 == _T_248) begin
                                      mem_51 <= _GEN_19;
                                    end else begin
                                      if (6'h33 == _T_243) begin
                                        mem_51 <= _GEN_18;
                                      end else begin
                                        if (6'h33 == _T_238) begin
                                          mem_51 <= _GEN_17;
                                        end else begin
                                          if (6'h33 == _T_233) begin
                                            mem_51 <= _GEN_16;
                                          end else begin
                                            if (6'h33 == _T_228) begin
                                              mem_51 <= _GEN_15;
                                            end else begin
                                              if (6'h33 == _T_223) begin
                                                mem_51 <= _GEN_14;
                                              end else begin
                                                if (6'h33 == _T_218) begin
                                                  mem_51 <= _GEN_13;
                                                end else begin
                                                  if (6'h33 == _T_213) begin
                                                    mem_51 <= _GEN_12;
                                                  end else begin
                                                    if (6'h33 == _T_208) begin
                                                      mem_51 <= _GEN_11;
                                                    end else begin
                                                      if (6'h33 == _T_203) begin
                                                        mem_51 <= _GEN_10;
                                                      end else begin
                                                        if (6'h33 == _T_198) begin
                                                          mem_51 <= _GEN_9;
                                                        end else begin
                                                          if (6'h33 == _T_193) begin
                                                            mem_51 <= _GEN_8;
                                                          end else begin
                                                            if (6'h33 == _T_188) begin
                                                              mem_51 <= _GEN_7;
                                                            end else begin
                                                              if (6'h33 == _T_183) begin
                                                                mem_51 <= _GEN_6;
                                                              end else begin
                                                                if (6'h33 == _T_178) begin
                                                                  mem_51 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h33 == _T_173) begin
                                                                    mem_51 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h33 == _T_168) begin
                                                                      mem_51 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h33 == _T_163) begin
                                                                        mem_51 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h33 == _T_158) begin
                                                                          mem_51 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h33 == _T_153) begin
                                                                            mem_51 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h33 == _T_308) begin
            mem_51 <= _GEN_31;
          end else begin
            if (6'h33 == _T_303) begin
              mem_51 <= _GEN_30;
            end else begin
              if (6'h33 == _T_298) begin
                mem_51 <= _GEN_29;
              end else begin
                if (6'h33 == _T_293) begin
                  mem_51 <= _GEN_28;
                end else begin
                  if (6'h33 == _T_288) begin
                    mem_51 <= _GEN_27;
                  end else begin
                    if (6'h33 == _T_283) begin
                      mem_51 <= _GEN_26;
                    end else begin
                      if (6'h33 == _T_278) begin
                        mem_51 <= _GEN_25;
                      end else begin
                        if (6'h33 == _T_273) begin
                          mem_51 <= _GEN_24;
                        end else begin
                          if (6'h33 == _T_268) begin
                            mem_51 <= _GEN_23;
                          end else begin
                            if (6'h33 == _T_263) begin
                              mem_51 <= _GEN_22;
                            end else begin
                              if (6'h33 == _T_258) begin
                                mem_51 <= _GEN_21;
                              end else begin
                                if (6'h33 == _T_253) begin
                                  mem_51 <= _GEN_20;
                                end else begin
                                  if (6'h33 == _T_248) begin
                                    mem_51 <= _GEN_19;
                                  end else begin
                                    if (6'h33 == _T_243) begin
                                      mem_51 <= _GEN_18;
                                    end else begin
                                      if (6'h33 == _T_238) begin
                                        mem_51 <= _GEN_17;
                                      end else begin
                                        if (6'h33 == _T_233) begin
                                          mem_51 <= _GEN_16;
                                        end else begin
                                          if (6'h33 == _T_228) begin
                                            mem_51 <= _GEN_15;
                                          end else begin
                                            if (6'h33 == _T_223) begin
                                              mem_51 <= _GEN_14;
                                            end else begin
                                              if (6'h33 == _T_218) begin
                                                mem_51 <= _GEN_13;
                                              end else begin
                                                if (6'h33 == _T_213) begin
                                                  mem_51 <= _GEN_12;
                                                end else begin
                                                  if (6'h33 == _T_208) begin
                                                    mem_51 <= _GEN_11;
                                                  end else begin
                                                    if (6'h33 == _T_203) begin
                                                      mem_51 <= _GEN_10;
                                                    end else begin
                                                      if (6'h33 == _T_198) begin
                                                        mem_51 <= _GEN_9;
                                                      end else begin
                                                        if (6'h33 == _T_193) begin
                                                          mem_51 <= _GEN_8;
                                                        end else begin
                                                          if (6'h33 == _T_188) begin
                                                            mem_51 <= _GEN_7;
                                                          end else begin
                                                            if (6'h33 == _T_183) begin
                                                              mem_51 <= _GEN_6;
                                                            end else begin
                                                              if (6'h33 == _T_178) begin
                                                                mem_51 <= _GEN_5;
                                                              end else begin
                                                                if (6'h33 == _T_173) begin
                                                                  mem_51 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h33 == _T_168) begin
                                                                    mem_51 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h33 == _T_163) begin
                                                                      mem_51 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h33 == _T_158) begin
                                                                        mem_51 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h33 == _T_153) begin
                                                                          mem_51 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h33 == _T_308) begin
          mem_51 <= _GEN_31;
        end else begin
          if (6'h33 == _T_303) begin
            mem_51 <= _GEN_30;
          end else begin
            if (6'h33 == _T_298) begin
              mem_51 <= _GEN_29;
            end else begin
              if (6'h33 == _T_293) begin
                mem_51 <= _GEN_28;
              end else begin
                if (6'h33 == _T_288) begin
                  mem_51 <= _GEN_27;
                end else begin
                  if (6'h33 == _T_283) begin
                    mem_51 <= _GEN_26;
                  end else begin
                    if (6'h33 == _T_278) begin
                      mem_51 <= _GEN_25;
                    end else begin
                      if (6'h33 == _T_273) begin
                        mem_51 <= _GEN_24;
                      end else begin
                        if (6'h33 == _T_268) begin
                          mem_51 <= _GEN_23;
                        end else begin
                          if (6'h33 == _T_263) begin
                            mem_51 <= _GEN_22;
                          end else begin
                            if (6'h33 == _T_258) begin
                              mem_51 <= _GEN_21;
                            end else begin
                              if (6'h33 == _T_253) begin
                                mem_51 <= _GEN_20;
                              end else begin
                                if (6'h33 == _T_248) begin
                                  mem_51 <= _GEN_19;
                                end else begin
                                  if (6'h33 == _T_243) begin
                                    mem_51 <= _GEN_18;
                                  end else begin
                                    if (6'h33 == _T_238) begin
                                      mem_51 <= _GEN_17;
                                    end else begin
                                      if (6'h33 == _T_233) begin
                                        mem_51 <= _GEN_16;
                                      end else begin
                                        if (6'h33 == _T_228) begin
                                          mem_51 <= _GEN_15;
                                        end else begin
                                          if (6'h33 == _T_223) begin
                                            mem_51 <= _GEN_14;
                                          end else begin
                                            if (6'h33 == _T_218) begin
                                              mem_51 <= _GEN_13;
                                            end else begin
                                              if (6'h33 == _T_213) begin
                                                mem_51 <= _GEN_12;
                                              end else begin
                                                if (6'h33 == _T_208) begin
                                                  mem_51 <= _GEN_11;
                                                end else begin
                                                  if (6'h33 == _T_203) begin
                                                    mem_51 <= _GEN_10;
                                                  end else begin
                                                    if (6'h33 == _T_198) begin
                                                      mem_51 <= _GEN_9;
                                                    end else begin
                                                      if (6'h33 == _T_193) begin
                                                        mem_51 <= _GEN_8;
                                                      end else begin
                                                        if (6'h33 == _T_188) begin
                                                          mem_51 <= _GEN_7;
                                                        end else begin
                                                          if (6'h33 == _T_183) begin
                                                            mem_51 <= _GEN_6;
                                                          end else begin
                                                            if (6'h33 == _T_178) begin
                                                              mem_51 <= _GEN_5;
                                                            end else begin
                                                              if (6'h33 == _T_173) begin
                                                                mem_51 <= _GEN_4;
                                                              end else begin
                                                                if (6'h33 == _T_168) begin
                                                                  mem_51 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h33 == _T_163) begin
                                                                    mem_51 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h33 == _T_158) begin
                                                                      mem_51 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h33 == _T_153) begin
                                                                        mem_51 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h34 == wPos) begin
            mem_52 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h34 == _T_308) begin
                mem_52 <= _GEN_31;
              end else begin
                if (6'h34 == _T_303) begin
                  mem_52 <= _GEN_30;
                end else begin
                  if (6'h34 == _T_298) begin
                    mem_52 <= _GEN_29;
                  end else begin
                    if (6'h34 == _T_293) begin
                      mem_52 <= _GEN_28;
                    end else begin
                      if (6'h34 == _T_288) begin
                        mem_52 <= _GEN_27;
                      end else begin
                        if (6'h34 == _T_283) begin
                          mem_52 <= _GEN_26;
                        end else begin
                          if (6'h34 == _T_278) begin
                            mem_52 <= _GEN_25;
                          end else begin
                            if (6'h34 == _T_273) begin
                              mem_52 <= _GEN_24;
                            end else begin
                              if (6'h34 == _T_268) begin
                                mem_52 <= _GEN_23;
                              end else begin
                                if (6'h34 == _T_263) begin
                                  mem_52 <= _GEN_22;
                                end else begin
                                  if (6'h34 == _T_258) begin
                                    mem_52 <= _GEN_21;
                                  end else begin
                                    if (6'h34 == _T_253) begin
                                      mem_52 <= _GEN_20;
                                    end else begin
                                      if (6'h34 == _T_248) begin
                                        mem_52 <= _GEN_19;
                                      end else begin
                                        if (6'h34 == _T_243) begin
                                          mem_52 <= _GEN_18;
                                        end else begin
                                          if (6'h34 == _T_238) begin
                                            mem_52 <= _GEN_17;
                                          end else begin
                                            if (6'h34 == _T_233) begin
                                              mem_52 <= _GEN_16;
                                            end else begin
                                              if (6'h34 == _T_228) begin
                                                mem_52 <= _GEN_15;
                                              end else begin
                                                if (6'h34 == _T_223) begin
                                                  mem_52 <= _GEN_14;
                                                end else begin
                                                  if (6'h34 == _T_218) begin
                                                    mem_52 <= _GEN_13;
                                                  end else begin
                                                    if (6'h34 == _T_213) begin
                                                      mem_52 <= _GEN_12;
                                                    end else begin
                                                      if (6'h34 == _T_208) begin
                                                        mem_52 <= _GEN_11;
                                                      end else begin
                                                        if (6'h34 == _T_203) begin
                                                          mem_52 <= _GEN_10;
                                                        end else begin
                                                          if (6'h34 == _T_198) begin
                                                            mem_52 <= _GEN_9;
                                                          end else begin
                                                            if (6'h34 == _T_193) begin
                                                              mem_52 <= _GEN_8;
                                                            end else begin
                                                              if (6'h34 == _T_188) begin
                                                                mem_52 <= _GEN_7;
                                                              end else begin
                                                                if (6'h34 == _T_183) begin
                                                                  mem_52 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h34 == _T_178) begin
                                                                    mem_52 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h34 == _T_173) begin
                                                                      mem_52 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h34 == _T_168) begin
                                                                        mem_52 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h34 == _T_163) begin
                                                                          mem_52 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h34 == _T_158) begin
                                                                            mem_52 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h34 == _T_153) begin
                                                                              mem_52 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h34 == _T_308) begin
              mem_52 <= _GEN_31;
            end else begin
              if (6'h34 == _T_303) begin
                mem_52 <= _GEN_30;
              end else begin
                if (6'h34 == _T_298) begin
                  mem_52 <= _GEN_29;
                end else begin
                  if (6'h34 == _T_293) begin
                    mem_52 <= _GEN_28;
                  end else begin
                    if (6'h34 == _T_288) begin
                      mem_52 <= _GEN_27;
                    end else begin
                      if (6'h34 == _T_283) begin
                        mem_52 <= _GEN_26;
                      end else begin
                        if (6'h34 == _T_278) begin
                          mem_52 <= _GEN_25;
                        end else begin
                          if (6'h34 == _T_273) begin
                            mem_52 <= _GEN_24;
                          end else begin
                            if (6'h34 == _T_268) begin
                              mem_52 <= _GEN_23;
                            end else begin
                              if (6'h34 == _T_263) begin
                                mem_52 <= _GEN_22;
                              end else begin
                                if (6'h34 == _T_258) begin
                                  mem_52 <= _GEN_21;
                                end else begin
                                  if (6'h34 == _T_253) begin
                                    mem_52 <= _GEN_20;
                                  end else begin
                                    if (6'h34 == _T_248) begin
                                      mem_52 <= _GEN_19;
                                    end else begin
                                      if (6'h34 == _T_243) begin
                                        mem_52 <= _GEN_18;
                                      end else begin
                                        if (6'h34 == _T_238) begin
                                          mem_52 <= _GEN_17;
                                        end else begin
                                          if (6'h34 == _T_233) begin
                                            mem_52 <= _GEN_16;
                                          end else begin
                                            if (6'h34 == _T_228) begin
                                              mem_52 <= _GEN_15;
                                            end else begin
                                              if (6'h34 == _T_223) begin
                                                mem_52 <= _GEN_14;
                                              end else begin
                                                if (6'h34 == _T_218) begin
                                                  mem_52 <= _GEN_13;
                                                end else begin
                                                  if (6'h34 == _T_213) begin
                                                    mem_52 <= _GEN_12;
                                                  end else begin
                                                    if (6'h34 == _T_208) begin
                                                      mem_52 <= _GEN_11;
                                                    end else begin
                                                      if (6'h34 == _T_203) begin
                                                        mem_52 <= _GEN_10;
                                                      end else begin
                                                        if (6'h34 == _T_198) begin
                                                          mem_52 <= _GEN_9;
                                                        end else begin
                                                          if (6'h34 == _T_193) begin
                                                            mem_52 <= _GEN_8;
                                                          end else begin
                                                            if (6'h34 == _T_188) begin
                                                              mem_52 <= _GEN_7;
                                                            end else begin
                                                              if (6'h34 == _T_183) begin
                                                                mem_52 <= _GEN_6;
                                                              end else begin
                                                                if (6'h34 == _T_178) begin
                                                                  mem_52 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h34 == _T_173) begin
                                                                    mem_52 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h34 == _T_168) begin
                                                                      mem_52 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h34 == _T_163) begin
                                                                        mem_52 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h34 == _T_158) begin
                                                                          mem_52 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h34 == _T_153) begin
                                                                            mem_52 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h34 == _T_308) begin
            mem_52 <= _GEN_31;
          end else begin
            if (6'h34 == _T_303) begin
              mem_52 <= _GEN_30;
            end else begin
              if (6'h34 == _T_298) begin
                mem_52 <= _GEN_29;
              end else begin
                if (6'h34 == _T_293) begin
                  mem_52 <= _GEN_28;
                end else begin
                  if (6'h34 == _T_288) begin
                    mem_52 <= _GEN_27;
                  end else begin
                    if (6'h34 == _T_283) begin
                      mem_52 <= _GEN_26;
                    end else begin
                      if (6'h34 == _T_278) begin
                        mem_52 <= _GEN_25;
                      end else begin
                        if (6'h34 == _T_273) begin
                          mem_52 <= _GEN_24;
                        end else begin
                          if (6'h34 == _T_268) begin
                            mem_52 <= _GEN_23;
                          end else begin
                            if (6'h34 == _T_263) begin
                              mem_52 <= _GEN_22;
                            end else begin
                              if (6'h34 == _T_258) begin
                                mem_52 <= _GEN_21;
                              end else begin
                                if (6'h34 == _T_253) begin
                                  mem_52 <= _GEN_20;
                                end else begin
                                  if (6'h34 == _T_248) begin
                                    mem_52 <= _GEN_19;
                                  end else begin
                                    if (6'h34 == _T_243) begin
                                      mem_52 <= _GEN_18;
                                    end else begin
                                      if (6'h34 == _T_238) begin
                                        mem_52 <= _GEN_17;
                                      end else begin
                                        if (6'h34 == _T_233) begin
                                          mem_52 <= _GEN_16;
                                        end else begin
                                          if (6'h34 == _T_228) begin
                                            mem_52 <= _GEN_15;
                                          end else begin
                                            if (6'h34 == _T_223) begin
                                              mem_52 <= _GEN_14;
                                            end else begin
                                              if (6'h34 == _T_218) begin
                                                mem_52 <= _GEN_13;
                                              end else begin
                                                if (6'h34 == _T_213) begin
                                                  mem_52 <= _GEN_12;
                                                end else begin
                                                  if (6'h34 == _T_208) begin
                                                    mem_52 <= _GEN_11;
                                                  end else begin
                                                    if (6'h34 == _T_203) begin
                                                      mem_52 <= _GEN_10;
                                                    end else begin
                                                      if (6'h34 == _T_198) begin
                                                        mem_52 <= _GEN_9;
                                                      end else begin
                                                        if (6'h34 == _T_193) begin
                                                          mem_52 <= _GEN_8;
                                                        end else begin
                                                          if (6'h34 == _T_188) begin
                                                            mem_52 <= _GEN_7;
                                                          end else begin
                                                            if (6'h34 == _T_183) begin
                                                              mem_52 <= _GEN_6;
                                                            end else begin
                                                              if (6'h34 == _T_178) begin
                                                                mem_52 <= _GEN_5;
                                                              end else begin
                                                                if (6'h34 == _T_173) begin
                                                                  mem_52 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h34 == _T_168) begin
                                                                    mem_52 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h34 == _T_163) begin
                                                                      mem_52 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h34 == _T_158) begin
                                                                        mem_52 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h34 == _T_153) begin
                                                                          mem_52 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h34 == _T_308) begin
          mem_52 <= _GEN_31;
        end else begin
          if (6'h34 == _T_303) begin
            mem_52 <= _GEN_30;
          end else begin
            if (6'h34 == _T_298) begin
              mem_52 <= _GEN_29;
            end else begin
              if (6'h34 == _T_293) begin
                mem_52 <= _GEN_28;
              end else begin
                if (6'h34 == _T_288) begin
                  mem_52 <= _GEN_27;
                end else begin
                  if (6'h34 == _T_283) begin
                    mem_52 <= _GEN_26;
                  end else begin
                    if (6'h34 == _T_278) begin
                      mem_52 <= _GEN_25;
                    end else begin
                      if (6'h34 == _T_273) begin
                        mem_52 <= _GEN_24;
                      end else begin
                        if (6'h34 == _T_268) begin
                          mem_52 <= _GEN_23;
                        end else begin
                          if (6'h34 == _T_263) begin
                            mem_52 <= _GEN_22;
                          end else begin
                            if (6'h34 == _T_258) begin
                              mem_52 <= _GEN_21;
                            end else begin
                              if (6'h34 == _T_253) begin
                                mem_52 <= _GEN_20;
                              end else begin
                                if (6'h34 == _T_248) begin
                                  mem_52 <= _GEN_19;
                                end else begin
                                  if (6'h34 == _T_243) begin
                                    mem_52 <= _GEN_18;
                                  end else begin
                                    if (6'h34 == _T_238) begin
                                      mem_52 <= _GEN_17;
                                    end else begin
                                      if (6'h34 == _T_233) begin
                                        mem_52 <= _GEN_16;
                                      end else begin
                                        if (6'h34 == _T_228) begin
                                          mem_52 <= _GEN_15;
                                        end else begin
                                          if (6'h34 == _T_223) begin
                                            mem_52 <= _GEN_14;
                                          end else begin
                                            if (6'h34 == _T_218) begin
                                              mem_52 <= _GEN_13;
                                            end else begin
                                              if (6'h34 == _T_213) begin
                                                mem_52 <= _GEN_12;
                                              end else begin
                                                if (6'h34 == _T_208) begin
                                                  mem_52 <= _GEN_11;
                                                end else begin
                                                  if (6'h34 == _T_203) begin
                                                    mem_52 <= _GEN_10;
                                                  end else begin
                                                    if (6'h34 == _T_198) begin
                                                      mem_52 <= _GEN_9;
                                                    end else begin
                                                      if (6'h34 == _T_193) begin
                                                        mem_52 <= _GEN_8;
                                                      end else begin
                                                        if (6'h34 == _T_188) begin
                                                          mem_52 <= _GEN_7;
                                                        end else begin
                                                          if (6'h34 == _T_183) begin
                                                            mem_52 <= _GEN_6;
                                                          end else begin
                                                            if (6'h34 == _T_178) begin
                                                              mem_52 <= _GEN_5;
                                                            end else begin
                                                              if (6'h34 == _T_173) begin
                                                                mem_52 <= _GEN_4;
                                                              end else begin
                                                                if (6'h34 == _T_168) begin
                                                                  mem_52 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h34 == _T_163) begin
                                                                    mem_52 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h34 == _T_158) begin
                                                                      mem_52 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h34 == _T_153) begin
                                                                        mem_52 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h35 == wPos) begin
            mem_53 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h35 == _T_308) begin
                mem_53 <= _GEN_31;
              end else begin
                if (6'h35 == _T_303) begin
                  mem_53 <= _GEN_30;
                end else begin
                  if (6'h35 == _T_298) begin
                    mem_53 <= _GEN_29;
                  end else begin
                    if (6'h35 == _T_293) begin
                      mem_53 <= _GEN_28;
                    end else begin
                      if (6'h35 == _T_288) begin
                        mem_53 <= _GEN_27;
                      end else begin
                        if (6'h35 == _T_283) begin
                          mem_53 <= _GEN_26;
                        end else begin
                          if (6'h35 == _T_278) begin
                            mem_53 <= _GEN_25;
                          end else begin
                            if (6'h35 == _T_273) begin
                              mem_53 <= _GEN_24;
                            end else begin
                              if (6'h35 == _T_268) begin
                                mem_53 <= _GEN_23;
                              end else begin
                                if (6'h35 == _T_263) begin
                                  mem_53 <= _GEN_22;
                                end else begin
                                  if (6'h35 == _T_258) begin
                                    mem_53 <= _GEN_21;
                                  end else begin
                                    if (6'h35 == _T_253) begin
                                      mem_53 <= _GEN_20;
                                    end else begin
                                      if (6'h35 == _T_248) begin
                                        mem_53 <= _GEN_19;
                                      end else begin
                                        if (6'h35 == _T_243) begin
                                          mem_53 <= _GEN_18;
                                        end else begin
                                          if (6'h35 == _T_238) begin
                                            mem_53 <= _GEN_17;
                                          end else begin
                                            if (6'h35 == _T_233) begin
                                              mem_53 <= _GEN_16;
                                            end else begin
                                              if (6'h35 == _T_228) begin
                                                mem_53 <= _GEN_15;
                                              end else begin
                                                if (6'h35 == _T_223) begin
                                                  mem_53 <= _GEN_14;
                                                end else begin
                                                  if (6'h35 == _T_218) begin
                                                    mem_53 <= _GEN_13;
                                                  end else begin
                                                    if (6'h35 == _T_213) begin
                                                      mem_53 <= _GEN_12;
                                                    end else begin
                                                      if (6'h35 == _T_208) begin
                                                        mem_53 <= _GEN_11;
                                                      end else begin
                                                        if (6'h35 == _T_203) begin
                                                          mem_53 <= _GEN_10;
                                                        end else begin
                                                          if (6'h35 == _T_198) begin
                                                            mem_53 <= _GEN_9;
                                                          end else begin
                                                            if (6'h35 == _T_193) begin
                                                              mem_53 <= _GEN_8;
                                                            end else begin
                                                              if (6'h35 == _T_188) begin
                                                                mem_53 <= _GEN_7;
                                                              end else begin
                                                                if (6'h35 == _T_183) begin
                                                                  mem_53 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h35 == _T_178) begin
                                                                    mem_53 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h35 == _T_173) begin
                                                                      mem_53 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h35 == _T_168) begin
                                                                        mem_53 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h35 == _T_163) begin
                                                                          mem_53 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h35 == _T_158) begin
                                                                            mem_53 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h35 == _T_153) begin
                                                                              mem_53 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h35 == _T_308) begin
              mem_53 <= _GEN_31;
            end else begin
              if (6'h35 == _T_303) begin
                mem_53 <= _GEN_30;
              end else begin
                if (6'h35 == _T_298) begin
                  mem_53 <= _GEN_29;
                end else begin
                  if (6'h35 == _T_293) begin
                    mem_53 <= _GEN_28;
                  end else begin
                    if (6'h35 == _T_288) begin
                      mem_53 <= _GEN_27;
                    end else begin
                      if (6'h35 == _T_283) begin
                        mem_53 <= _GEN_26;
                      end else begin
                        if (6'h35 == _T_278) begin
                          mem_53 <= _GEN_25;
                        end else begin
                          if (6'h35 == _T_273) begin
                            mem_53 <= _GEN_24;
                          end else begin
                            if (6'h35 == _T_268) begin
                              mem_53 <= _GEN_23;
                            end else begin
                              if (6'h35 == _T_263) begin
                                mem_53 <= _GEN_22;
                              end else begin
                                if (6'h35 == _T_258) begin
                                  mem_53 <= _GEN_21;
                                end else begin
                                  if (6'h35 == _T_253) begin
                                    mem_53 <= _GEN_20;
                                  end else begin
                                    if (6'h35 == _T_248) begin
                                      mem_53 <= _GEN_19;
                                    end else begin
                                      if (6'h35 == _T_243) begin
                                        mem_53 <= _GEN_18;
                                      end else begin
                                        if (6'h35 == _T_238) begin
                                          mem_53 <= _GEN_17;
                                        end else begin
                                          if (6'h35 == _T_233) begin
                                            mem_53 <= _GEN_16;
                                          end else begin
                                            if (6'h35 == _T_228) begin
                                              mem_53 <= _GEN_15;
                                            end else begin
                                              if (6'h35 == _T_223) begin
                                                mem_53 <= _GEN_14;
                                              end else begin
                                                if (6'h35 == _T_218) begin
                                                  mem_53 <= _GEN_13;
                                                end else begin
                                                  if (6'h35 == _T_213) begin
                                                    mem_53 <= _GEN_12;
                                                  end else begin
                                                    if (6'h35 == _T_208) begin
                                                      mem_53 <= _GEN_11;
                                                    end else begin
                                                      if (6'h35 == _T_203) begin
                                                        mem_53 <= _GEN_10;
                                                      end else begin
                                                        if (6'h35 == _T_198) begin
                                                          mem_53 <= _GEN_9;
                                                        end else begin
                                                          if (6'h35 == _T_193) begin
                                                            mem_53 <= _GEN_8;
                                                          end else begin
                                                            if (6'h35 == _T_188) begin
                                                              mem_53 <= _GEN_7;
                                                            end else begin
                                                              if (6'h35 == _T_183) begin
                                                                mem_53 <= _GEN_6;
                                                              end else begin
                                                                if (6'h35 == _T_178) begin
                                                                  mem_53 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h35 == _T_173) begin
                                                                    mem_53 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h35 == _T_168) begin
                                                                      mem_53 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h35 == _T_163) begin
                                                                        mem_53 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h35 == _T_158) begin
                                                                          mem_53 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h35 == _T_153) begin
                                                                            mem_53 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h35 == _T_308) begin
            mem_53 <= _GEN_31;
          end else begin
            if (6'h35 == _T_303) begin
              mem_53 <= _GEN_30;
            end else begin
              if (6'h35 == _T_298) begin
                mem_53 <= _GEN_29;
              end else begin
                if (6'h35 == _T_293) begin
                  mem_53 <= _GEN_28;
                end else begin
                  if (6'h35 == _T_288) begin
                    mem_53 <= _GEN_27;
                  end else begin
                    if (6'h35 == _T_283) begin
                      mem_53 <= _GEN_26;
                    end else begin
                      if (6'h35 == _T_278) begin
                        mem_53 <= _GEN_25;
                      end else begin
                        if (6'h35 == _T_273) begin
                          mem_53 <= _GEN_24;
                        end else begin
                          if (6'h35 == _T_268) begin
                            mem_53 <= _GEN_23;
                          end else begin
                            if (6'h35 == _T_263) begin
                              mem_53 <= _GEN_22;
                            end else begin
                              if (6'h35 == _T_258) begin
                                mem_53 <= _GEN_21;
                              end else begin
                                if (6'h35 == _T_253) begin
                                  mem_53 <= _GEN_20;
                                end else begin
                                  if (6'h35 == _T_248) begin
                                    mem_53 <= _GEN_19;
                                  end else begin
                                    if (6'h35 == _T_243) begin
                                      mem_53 <= _GEN_18;
                                    end else begin
                                      if (6'h35 == _T_238) begin
                                        mem_53 <= _GEN_17;
                                      end else begin
                                        if (6'h35 == _T_233) begin
                                          mem_53 <= _GEN_16;
                                        end else begin
                                          if (6'h35 == _T_228) begin
                                            mem_53 <= _GEN_15;
                                          end else begin
                                            if (6'h35 == _T_223) begin
                                              mem_53 <= _GEN_14;
                                            end else begin
                                              if (6'h35 == _T_218) begin
                                                mem_53 <= _GEN_13;
                                              end else begin
                                                if (6'h35 == _T_213) begin
                                                  mem_53 <= _GEN_12;
                                                end else begin
                                                  if (6'h35 == _T_208) begin
                                                    mem_53 <= _GEN_11;
                                                  end else begin
                                                    if (6'h35 == _T_203) begin
                                                      mem_53 <= _GEN_10;
                                                    end else begin
                                                      if (6'h35 == _T_198) begin
                                                        mem_53 <= _GEN_9;
                                                      end else begin
                                                        if (6'h35 == _T_193) begin
                                                          mem_53 <= _GEN_8;
                                                        end else begin
                                                          if (6'h35 == _T_188) begin
                                                            mem_53 <= _GEN_7;
                                                          end else begin
                                                            if (6'h35 == _T_183) begin
                                                              mem_53 <= _GEN_6;
                                                            end else begin
                                                              if (6'h35 == _T_178) begin
                                                                mem_53 <= _GEN_5;
                                                              end else begin
                                                                if (6'h35 == _T_173) begin
                                                                  mem_53 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h35 == _T_168) begin
                                                                    mem_53 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h35 == _T_163) begin
                                                                      mem_53 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h35 == _T_158) begin
                                                                        mem_53 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h35 == _T_153) begin
                                                                          mem_53 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h35 == _T_308) begin
          mem_53 <= _GEN_31;
        end else begin
          if (6'h35 == _T_303) begin
            mem_53 <= _GEN_30;
          end else begin
            if (6'h35 == _T_298) begin
              mem_53 <= _GEN_29;
            end else begin
              if (6'h35 == _T_293) begin
                mem_53 <= _GEN_28;
              end else begin
                if (6'h35 == _T_288) begin
                  mem_53 <= _GEN_27;
                end else begin
                  if (6'h35 == _T_283) begin
                    mem_53 <= _GEN_26;
                  end else begin
                    if (6'h35 == _T_278) begin
                      mem_53 <= _GEN_25;
                    end else begin
                      if (6'h35 == _T_273) begin
                        mem_53 <= _GEN_24;
                      end else begin
                        if (6'h35 == _T_268) begin
                          mem_53 <= _GEN_23;
                        end else begin
                          if (6'h35 == _T_263) begin
                            mem_53 <= _GEN_22;
                          end else begin
                            if (6'h35 == _T_258) begin
                              mem_53 <= _GEN_21;
                            end else begin
                              if (6'h35 == _T_253) begin
                                mem_53 <= _GEN_20;
                              end else begin
                                if (6'h35 == _T_248) begin
                                  mem_53 <= _GEN_19;
                                end else begin
                                  if (6'h35 == _T_243) begin
                                    mem_53 <= _GEN_18;
                                  end else begin
                                    if (6'h35 == _T_238) begin
                                      mem_53 <= _GEN_17;
                                    end else begin
                                      if (6'h35 == _T_233) begin
                                        mem_53 <= _GEN_16;
                                      end else begin
                                        if (6'h35 == _T_228) begin
                                          mem_53 <= _GEN_15;
                                        end else begin
                                          if (6'h35 == _T_223) begin
                                            mem_53 <= _GEN_14;
                                          end else begin
                                            if (6'h35 == _T_218) begin
                                              mem_53 <= _GEN_13;
                                            end else begin
                                              if (6'h35 == _T_213) begin
                                                mem_53 <= _GEN_12;
                                              end else begin
                                                if (6'h35 == _T_208) begin
                                                  mem_53 <= _GEN_11;
                                                end else begin
                                                  if (6'h35 == _T_203) begin
                                                    mem_53 <= _GEN_10;
                                                  end else begin
                                                    if (6'h35 == _T_198) begin
                                                      mem_53 <= _GEN_9;
                                                    end else begin
                                                      if (6'h35 == _T_193) begin
                                                        mem_53 <= _GEN_8;
                                                      end else begin
                                                        if (6'h35 == _T_188) begin
                                                          mem_53 <= _GEN_7;
                                                        end else begin
                                                          if (6'h35 == _T_183) begin
                                                            mem_53 <= _GEN_6;
                                                          end else begin
                                                            if (6'h35 == _T_178) begin
                                                              mem_53 <= _GEN_5;
                                                            end else begin
                                                              if (6'h35 == _T_173) begin
                                                                mem_53 <= _GEN_4;
                                                              end else begin
                                                                if (6'h35 == _T_168) begin
                                                                  mem_53 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h35 == _T_163) begin
                                                                    mem_53 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h35 == _T_158) begin
                                                                      mem_53 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h35 == _T_153) begin
                                                                        mem_53 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h36 == wPos) begin
            mem_54 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h36 == _T_308) begin
                mem_54 <= _GEN_31;
              end else begin
                if (6'h36 == _T_303) begin
                  mem_54 <= _GEN_30;
                end else begin
                  if (6'h36 == _T_298) begin
                    mem_54 <= _GEN_29;
                  end else begin
                    if (6'h36 == _T_293) begin
                      mem_54 <= _GEN_28;
                    end else begin
                      if (6'h36 == _T_288) begin
                        mem_54 <= _GEN_27;
                      end else begin
                        if (6'h36 == _T_283) begin
                          mem_54 <= _GEN_26;
                        end else begin
                          if (6'h36 == _T_278) begin
                            mem_54 <= _GEN_25;
                          end else begin
                            if (6'h36 == _T_273) begin
                              mem_54 <= _GEN_24;
                            end else begin
                              if (6'h36 == _T_268) begin
                                mem_54 <= _GEN_23;
                              end else begin
                                if (6'h36 == _T_263) begin
                                  mem_54 <= _GEN_22;
                                end else begin
                                  if (6'h36 == _T_258) begin
                                    mem_54 <= _GEN_21;
                                  end else begin
                                    if (6'h36 == _T_253) begin
                                      mem_54 <= _GEN_20;
                                    end else begin
                                      if (6'h36 == _T_248) begin
                                        mem_54 <= _GEN_19;
                                      end else begin
                                        if (6'h36 == _T_243) begin
                                          mem_54 <= _GEN_18;
                                        end else begin
                                          if (6'h36 == _T_238) begin
                                            mem_54 <= _GEN_17;
                                          end else begin
                                            if (6'h36 == _T_233) begin
                                              mem_54 <= _GEN_16;
                                            end else begin
                                              if (6'h36 == _T_228) begin
                                                mem_54 <= _GEN_15;
                                              end else begin
                                                if (6'h36 == _T_223) begin
                                                  mem_54 <= _GEN_14;
                                                end else begin
                                                  if (6'h36 == _T_218) begin
                                                    mem_54 <= _GEN_13;
                                                  end else begin
                                                    if (6'h36 == _T_213) begin
                                                      mem_54 <= _GEN_12;
                                                    end else begin
                                                      if (6'h36 == _T_208) begin
                                                        mem_54 <= _GEN_11;
                                                      end else begin
                                                        if (6'h36 == _T_203) begin
                                                          mem_54 <= _GEN_10;
                                                        end else begin
                                                          if (6'h36 == _T_198) begin
                                                            mem_54 <= _GEN_9;
                                                          end else begin
                                                            if (6'h36 == _T_193) begin
                                                              mem_54 <= _GEN_8;
                                                            end else begin
                                                              if (6'h36 == _T_188) begin
                                                                mem_54 <= _GEN_7;
                                                              end else begin
                                                                if (6'h36 == _T_183) begin
                                                                  mem_54 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h36 == _T_178) begin
                                                                    mem_54 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h36 == _T_173) begin
                                                                      mem_54 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h36 == _T_168) begin
                                                                        mem_54 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h36 == _T_163) begin
                                                                          mem_54 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h36 == _T_158) begin
                                                                            mem_54 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h36 == _T_153) begin
                                                                              mem_54 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h36 == _T_308) begin
              mem_54 <= _GEN_31;
            end else begin
              if (6'h36 == _T_303) begin
                mem_54 <= _GEN_30;
              end else begin
                if (6'h36 == _T_298) begin
                  mem_54 <= _GEN_29;
                end else begin
                  if (6'h36 == _T_293) begin
                    mem_54 <= _GEN_28;
                  end else begin
                    if (6'h36 == _T_288) begin
                      mem_54 <= _GEN_27;
                    end else begin
                      if (6'h36 == _T_283) begin
                        mem_54 <= _GEN_26;
                      end else begin
                        if (6'h36 == _T_278) begin
                          mem_54 <= _GEN_25;
                        end else begin
                          if (6'h36 == _T_273) begin
                            mem_54 <= _GEN_24;
                          end else begin
                            if (6'h36 == _T_268) begin
                              mem_54 <= _GEN_23;
                            end else begin
                              if (6'h36 == _T_263) begin
                                mem_54 <= _GEN_22;
                              end else begin
                                if (6'h36 == _T_258) begin
                                  mem_54 <= _GEN_21;
                                end else begin
                                  if (6'h36 == _T_253) begin
                                    mem_54 <= _GEN_20;
                                  end else begin
                                    if (6'h36 == _T_248) begin
                                      mem_54 <= _GEN_19;
                                    end else begin
                                      if (6'h36 == _T_243) begin
                                        mem_54 <= _GEN_18;
                                      end else begin
                                        if (6'h36 == _T_238) begin
                                          mem_54 <= _GEN_17;
                                        end else begin
                                          if (6'h36 == _T_233) begin
                                            mem_54 <= _GEN_16;
                                          end else begin
                                            if (6'h36 == _T_228) begin
                                              mem_54 <= _GEN_15;
                                            end else begin
                                              if (6'h36 == _T_223) begin
                                                mem_54 <= _GEN_14;
                                              end else begin
                                                if (6'h36 == _T_218) begin
                                                  mem_54 <= _GEN_13;
                                                end else begin
                                                  if (6'h36 == _T_213) begin
                                                    mem_54 <= _GEN_12;
                                                  end else begin
                                                    if (6'h36 == _T_208) begin
                                                      mem_54 <= _GEN_11;
                                                    end else begin
                                                      if (6'h36 == _T_203) begin
                                                        mem_54 <= _GEN_10;
                                                      end else begin
                                                        if (6'h36 == _T_198) begin
                                                          mem_54 <= _GEN_9;
                                                        end else begin
                                                          if (6'h36 == _T_193) begin
                                                            mem_54 <= _GEN_8;
                                                          end else begin
                                                            if (6'h36 == _T_188) begin
                                                              mem_54 <= _GEN_7;
                                                            end else begin
                                                              if (6'h36 == _T_183) begin
                                                                mem_54 <= _GEN_6;
                                                              end else begin
                                                                if (6'h36 == _T_178) begin
                                                                  mem_54 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h36 == _T_173) begin
                                                                    mem_54 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h36 == _T_168) begin
                                                                      mem_54 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h36 == _T_163) begin
                                                                        mem_54 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h36 == _T_158) begin
                                                                          mem_54 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h36 == _T_153) begin
                                                                            mem_54 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h36 == _T_308) begin
            mem_54 <= _GEN_31;
          end else begin
            if (6'h36 == _T_303) begin
              mem_54 <= _GEN_30;
            end else begin
              if (6'h36 == _T_298) begin
                mem_54 <= _GEN_29;
              end else begin
                if (6'h36 == _T_293) begin
                  mem_54 <= _GEN_28;
                end else begin
                  if (6'h36 == _T_288) begin
                    mem_54 <= _GEN_27;
                  end else begin
                    if (6'h36 == _T_283) begin
                      mem_54 <= _GEN_26;
                    end else begin
                      if (6'h36 == _T_278) begin
                        mem_54 <= _GEN_25;
                      end else begin
                        if (6'h36 == _T_273) begin
                          mem_54 <= _GEN_24;
                        end else begin
                          if (6'h36 == _T_268) begin
                            mem_54 <= _GEN_23;
                          end else begin
                            if (6'h36 == _T_263) begin
                              mem_54 <= _GEN_22;
                            end else begin
                              if (6'h36 == _T_258) begin
                                mem_54 <= _GEN_21;
                              end else begin
                                if (6'h36 == _T_253) begin
                                  mem_54 <= _GEN_20;
                                end else begin
                                  if (6'h36 == _T_248) begin
                                    mem_54 <= _GEN_19;
                                  end else begin
                                    if (6'h36 == _T_243) begin
                                      mem_54 <= _GEN_18;
                                    end else begin
                                      if (6'h36 == _T_238) begin
                                        mem_54 <= _GEN_17;
                                      end else begin
                                        if (6'h36 == _T_233) begin
                                          mem_54 <= _GEN_16;
                                        end else begin
                                          if (6'h36 == _T_228) begin
                                            mem_54 <= _GEN_15;
                                          end else begin
                                            if (6'h36 == _T_223) begin
                                              mem_54 <= _GEN_14;
                                            end else begin
                                              if (6'h36 == _T_218) begin
                                                mem_54 <= _GEN_13;
                                              end else begin
                                                if (6'h36 == _T_213) begin
                                                  mem_54 <= _GEN_12;
                                                end else begin
                                                  if (6'h36 == _T_208) begin
                                                    mem_54 <= _GEN_11;
                                                  end else begin
                                                    if (6'h36 == _T_203) begin
                                                      mem_54 <= _GEN_10;
                                                    end else begin
                                                      if (6'h36 == _T_198) begin
                                                        mem_54 <= _GEN_9;
                                                      end else begin
                                                        if (6'h36 == _T_193) begin
                                                          mem_54 <= _GEN_8;
                                                        end else begin
                                                          if (6'h36 == _T_188) begin
                                                            mem_54 <= _GEN_7;
                                                          end else begin
                                                            if (6'h36 == _T_183) begin
                                                              mem_54 <= _GEN_6;
                                                            end else begin
                                                              if (6'h36 == _T_178) begin
                                                                mem_54 <= _GEN_5;
                                                              end else begin
                                                                if (6'h36 == _T_173) begin
                                                                  mem_54 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h36 == _T_168) begin
                                                                    mem_54 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h36 == _T_163) begin
                                                                      mem_54 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h36 == _T_158) begin
                                                                        mem_54 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h36 == _T_153) begin
                                                                          mem_54 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h36 == _T_308) begin
          mem_54 <= _GEN_31;
        end else begin
          if (6'h36 == _T_303) begin
            mem_54 <= _GEN_30;
          end else begin
            if (6'h36 == _T_298) begin
              mem_54 <= _GEN_29;
            end else begin
              if (6'h36 == _T_293) begin
                mem_54 <= _GEN_28;
              end else begin
                if (6'h36 == _T_288) begin
                  mem_54 <= _GEN_27;
                end else begin
                  if (6'h36 == _T_283) begin
                    mem_54 <= _GEN_26;
                  end else begin
                    if (6'h36 == _T_278) begin
                      mem_54 <= _GEN_25;
                    end else begin
                      if (6'h36 == _T_273) begin
                        mem_54 <= _GEN_24;
                      end else begin
                        if (6'h36 == _T_268) begin
                          mem_54 <= _GEN_23;
                        end else begin
                          if (6'h36 == _T_263) begin
                            mem_54 <= _GEN_22;
                          end else begin
                            if (6'h36 == _T_258) begin
                              mem_54 <= _GEN_21;
                            end else begin
                              if (6'h36 == _T_253) begin
                                mem_54 <= _GEN_20;
                              end else begin
                                if (6'h36 == _T_248) begin
                                  mem_54 <= _GEN_19;
                                end else begin
                                  if (6'h36 == _T_243) begin
                                    mem_54 <= _GEN_18;
                                  end else begin
                                    if (6'h36 == _T_238) begin
                                      mem_54 <= _GEN_17;
                                    end else begin
                                      if (6'h36 == _T_233) begin
                                        mem_54 <= _GEN_16;
                                      end else begin
                                        if (6'h36 == _T_228) begin
                                          mem_54 <= _GEN_15;
                                        end else begin
                                          if (6'h36 == _T_223) begin
                                            mem_54 <= _GEN_14;
                                          end else begin
                                            if (6'h36 == _T_218) begin
                                              mem_54 <= _GEN_13;
                                            end else begin
                                              if (6'h36 == _T_213) begin
                                                mem_54 <= _GEN_12;
                                              end else begin
                                                if (6'h36 == _T_208) begin
                                                  mem_54 <= _GEN_11;
                                                end else begin
                                                  if (6'h36 == _T_203) begin
                                                    mem_54 <= _GEN_10;
                                                  end else begin
                                                    if (6'h36 == _T_198) begin
                                                      mem_54 <= _GEN_9;
                                                    end else begin
                                                      if (6'h36 == _T_193) begin
                                                        mem_54 <= _GEN_8;
                                                      end else begin
                                                        if (6'h36 == _T_188) begin
                                                          mem_54 <= _GEN_7;
                                                        end else begin
                                                          if (6'h36 == _T_183) begin
                                                            mem_54 <= _GEN_6;
                                                          end else begin
                                                            if (6'h36 == _T_178) begin
                                                              mem_54 <= _GEN_5;
                                                            end else begin
                                                              if (6'h36 == _T_173) begin
                                                                mem_54 <= _GEN_4;
                                                              end else begin
                                                                if (6'h36 == _T_168) begin
                                                                  mem_54 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h36 == _T_163) begin
                                                                    mem_54 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h36 == _T_158) begin
                                                                      mem_54 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h36 == _T_153) begin
                                                                        mem_54 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h37 == wPos) begin
            mem_55 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h37 == _T_308) begin
                mem_55 <= _GEN_31;
              end else begin
                if (6'h37 == _T_303) begin
                  mem_55 <= _GEN_30;
                end else begin
                  if (6'h37 == _T_298) begin
                    mem_55 <= _GEN_29;
                  end else begin
                    if (6'h37 == _T_293) begin
                      mem_55 <= _GEN_28;
                    end else begin
                      if (6'h37 == _T_288) begin
                        mem_55 <= _GEN_27;
                      end else begin
                        if (6'h37 == _T_283) begin
                          mem_55 <= _GEN_26;
                        end else begin
                          if (6'h37 == _T_278) begin
                            mem_55 <= _GEN_25;
                          end else begin
                            if (6'h37 == _T_273) begin
                              mem_55 <= _GEN_24;
                            end else begin
                              if (6'h37 == _T_268) begin
                                mem_55 <= _GEN_23;
                              end else begin
                                if (6'h37 == _T_263) begin
                                  mem_55 <= _GEN_22;
                                end else begin
                                  if (6'h37 == _T_258) begin
                                    mem_55 <= _GEN_21;
                                  end else begin
                                    if (6'h37 == _T_253) begin
                                      mem_55 <= _GEN_20;
                                    end else begin
                                      if (6'h37 == _T_248) begin
                                        mem_55 <= _GEN_19;
                                      end else begin
                                        if (6'h37 == _T_243) begin
                                          mem_55 <= _GEN_18;
                                        end else begin
                                          if (6'h37 == _T_238) begin
                                            mem_55 <= _GEN_17;
                                          end else begin
                                            if (6'h37 == _T_233) begin
                                              mem_55 <= _GEN_16;
                                            end else begin
                                              if (6'h37 == _T_228) begin
                                                mem_55 <= _GEN_15;
                                              end else begin
                                                if (6'h37 == _T_223) begin
                                                  mem_55 <= _GEN_14;
                                                end else begin
                                                  if (6'h37 == _T_218) begin
                                                    mem_55 <= _GEN_13;
                                                  end else begin
                                                    if (6'h37 == _T_213) begin
                                                      mem_55 <= _GEN_12;
                                                    end else begin
                                                      if (6'h37 == _T_208) begin
                                                        mem_55 <= _GEN_11;
                                                      end else begin
                                                        if (6'h37 == _T_203) begin
                                                          mem_55 <= _GEN_10;
                                                        end else begin
                                                          if (6'h37 == _T_198) begin
                                                            mem_55 <= _GEN_9;
                                                          end else begin
                                                            if (6'h37 == _T_193) begin
                                                              mem_55 <= _GEN_8;
                                                            end else begin
                                                              if (6'h37 == _T_188) begin
                                                                mem_55 <= _GEN_7;
                                                              end else begin
                                                                if (6'h37 == _T_183) begin
                                                                  mem_55 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h37 == _T_178) begin
                                                                    mem_55 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h37 == _T_173) begin
                                                                      mem_55 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h37 == _T_168) begin
                                                                        mem_55 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h37 == _T_163) begin
                                                                          mem_55 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h37 == _T_158) begin
                                                                            mem_55 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h37 == _T_153) begin
                                                                              mem_55 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h37 == _T_308) begin
              mem_55 <= _GEN_31;
            end else begin
              if (6'h37 == _T_303) begin
                mem_55 <= _GEN_30;
              end else begin
                if (6'h37 == _T_298) begin
                  mem_55 <= _GEN_29;
                end else begin
                  if (6'h37 == _T_293) begin
                    mem_55 <= _GEN_28;
                  end else begin
                    if (6'h37 == _T_288) begin
                      mem_55 <= _GEN_27;
                    end else begin
                      if (6'h37 == _T_283) begin
                        mem_55 <= _GEN_26;
                      end else begin
                        if (6'h37 == _T_278) begin
                          mem_55 <= _GEN_25;
                        end else begin
                          if (6'h37 == _T_273) begin
                            mem_55 <= _GEN_24;
                          end else begin
                            if (6'h37 == _T_268) begin
                              mem_55 <= _GEN_23;
                            end else begin
                              if (6'h37 == _T_263) begin
                                mem_55 <= _GEN_22;
                              end else begin
                                if (6'h37 == _T_258) begin
                                  mem_55 <= _GEN_21;
                                end else begin
                                  if (6'h37 == _T_253) begin
                                    mem_55 <= _GEN_20;
                                  end else begin
                                    if (6'h37 == _T_248) begin
                                      mem_55 <= _GEN_19;
                                    end else begin
                                      if (6'h37 == _T_243) begin
                                        mem_55 <= _GEN_18;
                                      end else begin
                                        if (6'h37 == _T_238) begin
                                          mem_55 <= _GEN_17;
                                        end else begin
                                          if (6'h37 == _T_233) begin
                                            mem_55 <= _GEN_16;
                                          end else begin
                                            if (6'h37 == _T_228) begin
                                              mem_55 <= _GEN_15;
                                            end else begin
                                              if (6'h37 == _T_223) begin
                                                mem_55 <= _GEN_14;
                                              end else begin
                                                if (6'h37 == _T_218) begin
                                                  mem_55 <= _GEN_13;
                                                end else begin
                                                  if (6'h37 == _T_213) begin
                                                    mem_55 <= _GEN_12;
                                                  end else begin
                                                    if (6'h37 == _T_208) begin
                                                      mem_55 <= _GEN_11;
                                                    end else begin
                                                      if (6'h37 == _T_203) begin
                                                        mem_55 <= _GEN_10;
                                                      end else begin
                                                        if (6'h37 == _T_198) begin
                                                          mem_55 <= _GEN_9;
                                                        end else begin
                                                          if (6'h37 == _T_193) begin
                                                            mem_55 <= _GEN_8;
                                                          end else begin
                                                            if (6'h37 == _T_188) begin
                                                              mem_55 <= _GEN_7;
                                                            end else begin
                                                              if (6'h37 == _T_183) begin
                                                                mem_55 <= _GEN_6;
                                                              end else begin
                                                                if (6'h37 == _T_178) begin
                                                                  mem_55 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h37 == _T_173) begin
                                                                    mem_55 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h37 == _T_168) begin
                                                                      mem_55 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h37 == _T_163) begin
                                                                        mem_55 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h37 == _T_158) begin
                                                                          mem_55 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h37 == _T_153) begin
                                                                            mem_55 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h37 == _T_308) begin
            mem_55 <= _GEN_31;
          end else begin
            if (6'h37 == _T_303) begin
              mem_55 <= _GEN_30;
            end else begin
              if (6'h37 == _T_298) begin
                mem_55 <= _GEN_29;
              end else begin
                if (6'h37 == _T_293) begin
                  mem_55 <= _GEN_28;
                end else begin
                  if (6'h37 == _T_288) begin
                    mem_55 <= _GEN_27;
                  end else begin
                    if (6'h37 == _T_283) begin
                      mem_55 <= _GEN_26;
                    end else begin
                      if (6'h37 == _T_278) begin
                        mem_55 <= _GEN_25;
                      end else begin
                        if (6'h37 == _T_273) begin
                          mem_55 <= _GEN_24;
                        end else begin
                          if (6'h37 == _T_268) begin
                            mem_55 <= _GEN_23;
                          end else begin
                            if (6'h37 == _T_263) begin
                              mem_55 <= _GEN_22;
                            end else begin
                              if (6'h37 == _T_258) begin
                                mem_55 <= _GEN_21;
                              end else begin
                                if (6'h37 == _T_253) begin
                                  mem_55 <= _GEN_20;
                                end else begin
                                  if (6'h37 == _T_248) begin
                                    mem_55 <= _GEN_19;
                                  end else begin
                                    if (6'h37 == _T_243) begin
                                      mem_55 <= _GEN_18;
                                    end else begin
                                      if (6'h37 == _T_238) begin
                                        mem_55 <= _GEN_17;
                                      end else begin
                                        if (6'h37 == _T_233) begin
                                          mem_55 <= _GEN_16;
                                        end else begin
                                          if (6'h37 == _T_228) begin
                                            mem_55 <= _GEN_15;
                                          end else begin
                                            if (6'h37 == _T_223) begin
                                              mem_55 <= _GEN_14;
                                            end else begin
                                              if (6'h37 == _T_218) begin
                                                mem_55 <= _GEN_13;
                                              end else begin
                                                if (6'h37 == _T_213) begin
                                                  mem_55 <= _GEN_12;
                                                end else begin
                                                  if (6'h37 == _T_208) begin
                                                    mem_55 <= _GEN_11;
                                                  end else begin
                                                    if (6'h37 == _T_203) begin
                                                      mem_55 <= _GEN_10;
                                                    end else begin
                                                      if (6'h37 == _T_198) begin
                                                        mem_55 <= _GEN_9;
                                                      end else begin
                                                        if (6'h37 == _T_193) begin
                                                          mem_55 <= _GEN_8;
                                                        end else begin
                                                          if (6'h37 == _T_188) begin
                                                            mem_55 <= _GEN_7;
                                                          end else begin
                                                            if (6'h37 == _T_183) begin
                                                              mem_55 <= _GEN_6;
                                                            end else begin
                                                              if (6'h37 == _T_178) begin
                                                                mem_55 <= _GEN_5;
                                                              end else begin
                                                                if (6'h37 == _T_173) begin
                                                                  mem_55 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h37 == _T_168) begin
                                                                    mem_55 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h37 == _T_163) begin
                                                                      mem_55 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h37 == _T_158) begin
                                                                        mem_55 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h37 == _T_153) begin
                                                                          mem_55 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h37 == _T_308) begin
          mem_55 <= _GEN_31;
        end else begin
          if (6'h37 == _T_303) begin
            mem_55 <= _GEN_30;
          end else begin
            if (6'h37 == _T_298) begin
              mem_55 <= _GEN_29;
            end else begin
              if (6'h37 == _T_293) begin
                mem_55 <= _GEN_28;
              end else begin
                if (6'h37 == _T_288) begin
                  mem_55 <= _GEN_27;
                end else begin
                  if (6'h37 == _T_283) begin
                    mem_55 <= _GEN_26;
                  end else begin
                    if (6'h37 == _T_278) begin
                      mem_55 <= _GEN_25;
                    end else begin
                      if (6'h37 == _T_273) begin
                        mem_55 <= _GEN_24;
                      end else begin
                        if (6'h37 == _T_268) begin
                          mem_55 <= _GEN_23;
                        end else begin
                          if (6'h37 == _T_263) begin
                            mem_55 <= _GEN_22;
                          end else begin
                            if (6'h37 == _T_258) begin
                              mem_55 <= _GEN_21;
                            end else begin
                              if (6'h37 == _T_253) begin
                                mem_55 <= _GEN_20;
                              end else begin
                                if (6'h37 == _T_248) begin
                                  mem_55 <= _GEN_19;
                                end else begin
                                  if (6'h37 == _T_243) begin
                                    mem_55 <= _GEN_18;
                                  end else begin
                                    if (6'h37 == _T_238) begin
                                      mem_55 <= _GEN_17;
                                    end else begin
                                      if (6'h37 == _T_233) begin
                                        mem_55 <= _GEN_16;
                                      end else begin
                                        if (6'h37 == _T_228) begin
                                          mem_55 <= _GEN_15;
                                        end else begin
                                          if (6'h37 == _T_223) begin
                                            mem_55 <= _GEN_14;
                                          end else begin
                                            if (6'h37 == _T_218) begin
                                              mem_55 <= _GEN_13;
                                            end else begin
                                              if (6'h37 == _T_213) begin
                                                mem_55 <= _GEN_12;
                                              end else begin
                                                if (6'h37 == _T_208) begin
                                                  mem_55 <= _GEN_11;
                                                end else begin
                                                  if (6'h37 == _T_203) begin
                                                    mem_55 <= _GEN_10;
                                                  end else begin
                                                    if (6'h37 == _T_198) begin
                                                      mem_55 <= _GEN_9;
                                                    end else begin
                                                      if (6'h37 == _T_193) begin
                                                        mem_55 <= _GEN_8;
                                                      end else begin
                                                        if (6'h37 == _T_188) begin
                                                          mem_55 <= _GEN_7;
                                                        end else begin
                                                          if (6'h37 == _T_183) begin
                                                            mem_55 <= _GEN_6;
                                                          end else begin
                                                            if (6'h37 == _T_178) begin
                                                              mem_55 <= _GEN_5;
                                                            end else begin
                                                              if (6'h37 == _T_173) begin
                                                                mem_55 <= _GEN_4;
                                                              end else begin
                                                                if (6'h37 == _T_168) begin
                                                                  mem_55 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h37 == _T_163) begin
                                                                    mem_55 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h37 == _T_158) begin
                                                                      mem_55 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h37 == _T_153) begin
                                                                        mem_55 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h38 == wPos) begin
            mem_56 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h38 == _T_308) begin
                mem_56 <= _GEN_31;
              end else begin
                if (6'h38 == _T_303) begin
                  mem_56 <= _GEN_30;
                end else begin
                  if (6'h38 == _T_298) begin
                    mem_56 <= _GEN_29;
                  end else begin
                    if (6'h38 == _T_293) begin
                      mem_56 <= _GEN_28;
                    end else begin
                      if (6'h38 == _T_288) begin
                        mem_56 <= _GEN_27;
                      end else begin
                        if (6'h38 == _T_283) begin
                          mem_56 <= _GEN_26;
                        end else begin
                          if (6'h38 == _T_278) begin
                            mem_56 <= _GEN_25;
                          end else begin
                            if (6'h38 == _T_273) begin
                              mem_56 <= _GEN_24;
                            end else begin
                              if (6'h38 == _T_268) begin
                                mem_56 <= _GEN_23;
                              end else begin
                                if (6'h38 == _T_263) begin
                                  mem_56 <= _GEN_22;
                                end else begin
                                  if (6'h38 == _T_258) begin
                                    mem_56 <= _GEN_21;
                                  end else begin
                                    if (6'h38 == _T_253) begin
                                      mem_56 <= _GEN_20;
                                    end else begin
                                      if (6'h38 == _T_248) begin
                                        mem_56 <= _GEN_19;
                                      end else begin
                                        if (6'h38 == _T_243) begin
                                          mem_56 <= _GEN_18;
                                        end else begin
                                          if (6'h38 == _T_238) begin
                                            mem_56 <= _GEN_17;
                                          end else begin
                                            if (6'h38 == _T_233) begin
                                              mem_56 <= _GEN_16;
                                            end else begin
                                              if (6'h38 == _T_228) begin
                                                mem_56 <= _GEN_15;
                                              end else begin
                                                if (6'h38 == _T_223) begin
                                                  mem_56 <= _GEN_14;
                                                end else begin
                                                  if (6'h38 == _T_218) begin
                                                    mem_56 <= _GEN_13;
                                                  end else begin
                                                    if (6'h38 == _T_213) begin
                                                      mem_56 <= _GEN_12;
                                                    end else begin
                                                      if (6'h38 == _T_208) begin
                                                        mem_56 <= _GEN_11;
                                                      end else begin
                                                        if (6'h38 == _T_203) begin
                                                          mem_56 <= _GEN_10;
                                                        end else begin
                                                          if (6'h38 == _T_198) begin
                                                            mem_56 <= _GEN_9;
                                                          end else begin
                                                            if (6'h38 == _T_193) begin
                                                              mem_56 <= _GEN_8;
                                                            end else begin
                                                              if (6'h38 == _T_188) begin
                                                                mem_56 <= _GEN_7;
                                                              end else begin
                                                                if (6'h38 == _T_183) begin
                                                                  mem_56 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h38 == _T_178) begin
                                                                    mem_56 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h38 == _T_173) begin
                                                                      mem_56 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h38 == _T_168) begin
                                                                        mem_56 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h38 == _T_163) begin
                                                                          mem_56 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h38 == _T_158) begin
                                                                            mem_56 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h38 == _T_153) begin
                                                                              mem_56 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h38 == _T_308) begin
              mem_56 <= _GEN_31;
            end else begin
              if (6'h38 == _T_303) begin
                mem_56 <= _GEN_30;
              end else begin
                if (6'h38 == _T_298) begin
                  mem_56 <= _GEN_29;
                end else begin
                  if (6'h38 == _T_293) begin
                    mem_56 <= _GEN_28;
                  end else begin
                    if (6'h38 == _T_288) begin
                      mem_56 <= _GEN_27;
                    end else begin
                      if (6'h38 == _T_283) begin
                        mem_56 <= _GEN_26;
                      end else begin
                        if (6'h38 == _T_278) begin
                          mem_56 <= _GEN_25;
                        end else begin
                          if (6'h38 == _T_273) begin
                            mem_56 <= _GEN_24;
                          end else begin
                            if (6'h38 == _T_268) begin
                              mem_56 <= _GEN_23;
                            end else begin
                              if (6'h38 == _T_263) begin
                                mem_56 <= _GEN_22;
                              end else begin
                                if (6'h38 == _T_258) begin
                                  mem_56 <= _GEN_21;
                                end else begin
                                  if (6'h38 == _T_253) begin
                                    mem_56 <= _GEN_20;
                                  end else begin
                                    if (6'h38 == _T_248) begin
                                      mem_56 <= _GEN_19;
                                    end else begin
                                      if (6'h38 == _T_243) begin
                                        mem_56 <= _GEN_18;
                                      end else begin
                                        if (6'h38 == _T_238) begin
                                          mem_56 <= _GEN_17;
                                        end else begin
                                          if (6'h38 == _T_233) begin
                                            mem_56 <= _GEN_16;
                                          end else begin
                                            if (6'h38 == _T_228) begin
                                              mem_56 <= _GEN_15;
                                            end else begin
                                              if (6'h38 == _T_223) begin
                                                mem_56 <= _GEN_14;
                                              end else begin
                                                if (6'h38 == _T_218) begin
                                                  mem_56 <= _GEN_13;
                                                end else begin
                                                  if (6'h38 == _T_213) begin
                                                    mem_56 <= _GEN_12;
                                                  end else begin
                                                    if (6'h38 == _T_208) begin
                                                      mem_56 <= _GEN_11;
                                                    end else begin
                                                      if (6'h38 == _T_203) begin
                                                        mem_56 <= _GEN_10;
                                                      end else begin
                                                        if (6'h38 == _T_198) begin
                                                          mem_56 <= _GEN_9;
                                                        end else begin
                                                          if (6'h38 == _T_193) begin
                                                            mem_56 <= _GEN_8;
                                                          end else begin
                                                            if (6'h38 == _T_188) begin
                                                              mem_56 <= _GEN_7;
                                                            end else begin
                                                              if (6'h38 == _T_183) begin
                                                                mem_56 <= _GEN_6;
                                                              end else begin
                                                                if (6'h38 == _T_178) begin
                                                                  mem_56 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h38 == _T_173) begin
                                                                    mem_56 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h38 == _T_168) begin
                                                                      mem_56 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h38 == _T_163) begin
                                                                        mem_56 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h38 == _T_158) begin
                                                                          mem_56 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h38 == _T_153) begin
                                                                            mem_56 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h38 == _T_308) begin
            mem_56 <= _GEN_31;
          end else begin
            if (6'h38 == _T_303) begin
              mem_56 <= _GEN_30;
            end else begin
              if (6'h38 == _T_298) begin
                mem_56 <= _GEN_29;
              end else begin
                if (6'h38 == _T_293) begin
                  mem_56 <= _GEN_28;
                end else begin
                  if (6'h38 == _T_288) begin
                    mem_56 <= _GEN_27;
                  end else begin
                    if (6'h38 == _T_283) begin
                      mem_56 <= _GEN_26;
                    end else begin
                      if (6'h38 == _T_278) begin
                        mem_56 <= _GEN_25;
                      end else begin
                        if (6'h38 == _T_273) begin
                          mem_56 <= _GEN_24;
                        end else begin
                          if (6'h38 == _T_268) begin
                            mem_56 <= _GEN_23;
                          end else begin
                            if (6'h38 == _T_263) begin
                              mem_56 <= _GEN_22;
                            end else begin
                              if (6'h38 == _T_258) begin
                                mem_56 <= _GEN_21;
                              end else begin
                                if (6'h38 == _T_253) begin
                                  mem_56 <= _GEN_20;
                                end else begin
                                  if (6'h38 == _T_248) begin
                                    mem_56 <= _GEN_19;
                                  end else begin
                                    if (6'h38 == _T_243) begin
                                      mem_56 <= _GEN_18;
                                    end else begin
                                      if (6'h38 == _T_238) begin
                                        mem_56 <= _GEN_17;
                                      end else begin
                                        if (6'h38 == _T_233) begin
                                          mem_56 <= _GEN_16;
                                        end else begin
                                          if (6'h38 == _T_228) begin
                                            mem_56 <= _GEN_15;
                                          end else begin
                                            if (6'h38 == _T_223) begin
                                              mem_56 <= _GEN_14;
                                            end else begin
                                              if (6'h38 == _T_218) begin
                                                mem_56 <= _GEN_13;
                                              end else begin
                                                if (6'h38 == _T_213) begin
                                                  mem_56 <= _GEN_12;
                                                end else begin
                                                  if (6'h38 == _T_208) begin
                                                    mem_56 <= _GEN_11;
                                                  end else begin
                                                    if (6'h38 == _T_203) begin
                                                      mem_56 <= _GEN_10;
                                                    end else begin
                                                      if (6'h38 == _T_198) begin
                                                        mem_56 <= _GEN_9;
                                                      end else begin
                                                        if (6'h38 == _T_193) begin
                                                          mem_56 <= _GEN_8;
                                                        end else begin
                                                          if (6'h38 == _T_188) begin
                                                            mem_56 <= _GEN_7;
                                                          end else begin
                                                            if (6'h38 == _T_183) begin
                                                              mem_56 <= _GEN_6;
                                                            end else begin
                                                              if (6'h38 == _T_178) begin
                                                                mem_56 <= _GEN_5;
                                                              end else begin
                                                                if (6'h38 == _T_173) begin
                                                                  mem_56 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h38 == _T_168) begin
                                                                    mem_56 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h38 == _T_163) begin
                                                                      mem_56 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h38 == _T_158) begin
                                                                        mem_56 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h38 == _T_153) begin
                                                                          mem_56 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h38 == _T_308) begin
          mem_56 <= _GEN_31;
        end else begin
          if (6'h38 == _T_303) begin
            mem_56 <= _GEN_30;
          end else begin
            if (6'h38 == _T_298) begin
              mem_56 <= _GEN_29;
            end else begin
              if (6'h38 == _T_293) begin
                mem_56 <= _GEN_28;
              end else begin
                if (6'h38 == _T_288) begin
                  mem_56 <= _GEN_27;
                end else begin
                  if (6'h38 == _T_283) begin
                    mem_56 <= _GEN_26;
                  end else begin
                    if (6'h38 == _T_278) begin
                      mem_56 <= _GEN_25;
                    end else begin
                      if (6'h38 == _T_273) begin
                        mem_56 <= _GEN_24;
                      end else begin
                        if (6'h38 == _T_268) begin
                          mem_56 <= _GEN_23;
                        end else begin
                          if (6'h38 == _T_263) begin
                            mem_56 <= _GEN_22;
                          end else begin
                            if (6'h38 == _T_258) begin
                              mem_56 <= _GEN_21;
                            end else begin
                              if (6'h38 == _T_253) begin
                                mem_56 <= _GEN_20;
                              end else begin
                                if (6'h38 == _T_248) begin
                                  mem_56 <= _GEN_19;
                                end else begin
                                  if (6'h38 == _T_243) begin
                                    mem_56 <= _GEN_18;
                                  end else begin
                                    if (6'h38 == _T_238) begin
                                      mem_56 <= _GEN_17;
                                    end else begin
                                      if (6'h38 == _T_233) begin
                                        mem_56 <= _GEN_16;
                                      end else begin
                                        if (6'h38 == _T_228) begin
                                          mem_56 <= _GEN_15;
                                        end else begin
                                          if (6'h38 == _T_223) begin
                                            mem_56 <= _GEN_14;
                                          end else begin
                                            if (6'h38 == _T_218) begin
                                              mem_56 <= _GEN_13;
                                            end else begin
                                              if (6'h38 == _T_213) begin
                                                mem_56 <= _GEN_12;
                                              end else begin
                                                if (6'h38 == _T_208) begin
                                                  mem_56 <= _GEN_11;
                                                end else begin
                                                  if (6'h38 == _T_203) begin
                                                    mem_56 <= _GEN_10;
                                                  end else begin
                                                    if (6'h38 == _T_198) begin
                                                      mem_56 <= _GEN_9;
                                                    end else begin
                                                      if (6'h38 == _T_193) begin
                                                        mem_56 <= _GEN_8;
                                                      end else begin
                                                        if (6'h38 == _T_188) begin
                                                          mem_56 <= _GEN_7;
                                                        end else begin
                                                          if (6'h38 == _T_183) begin
                                                            mem_56 <= _GEN_6;
                                                          end else begin
                                                            if (6'h38 == _T_178) begin
                                                              mem_56 <= _GEN_5;
                                                            end else begin
                                                              if (6'h38 == _T_173) begin
                                                                mem_56 <= _GEN_4;
                                                              end else begin
                                                                if (6'h38 == _T_168) begin
                                                                  mem_56 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h38 == _T_163) begin
                                                                    mem_56 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h38 == _T_158) begin
                                                                      mem_56 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h38 == _T_153) begin
                                                                        mem_56 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h39 == wPos) begin
            mem_57 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h39 == _T_308) begin
                mem_57 <= _GEN_31;
              end else begin
                if (6'h39 == _T_303) begin
                  mem_57 <= _GEN_30;
                end else begin
                  if (6'h39 == _T_298) begin
                    mem_57 <= _GEN_29;
                  end else begin
                    if (6'h39 == _T_293) begin
                      mem_57 <= _GEN_28;
                    end else begin
                      if (6'h39 == _T_288) begin
                        mem_57 <= _GEN_27;
                      end else begin
                        if (6'h39 == _T_283) begin
                          mem_57 <= _GEN_26;
                        end else begin
                          if (6'h39 == _T_278) begin
                            mem_57 <= _GEN_25;
                          end else begin
                            if (6'h39 == _T_273) begin
                              mem_57 <= _GEN_24;
                            end else begin
                              if (6'h39 == _T_268) begin
                                mem_57 <= _GEN_23;
                              end else begin
                                if (6'h39 == _T_263) begin
                                  mem_57 <= _GEN_22;
                                end else begin
                                  if (6'h39 == _T_258) begin
                                    mem_57 <= _GEN_21;
                                  end else begin
                                    if (6'h39 == _T_253) begin
                                      mem_57 <= _GEN_20;
                                    end else begin
                                      if (6'h39 == _T_248) begin
                                        mem_57 <= _GEN_19;
                                      end else begin
                                        if (6'h39 == _T_243) begin
                                          mem_57 <= _GEN_18;
                                        end else begin
                                          if (6'h39 == _T_238) begin
                                            mem_57 <= _GEN_17;
                                          end else begin
                                            if (6'h39 == _T_233) begin
                                              mem_57 <= _GEN_16;
                                            end else begin
                                              if (6'h39 == _T_228) begin
                                                mem_57 <= _GEN_15;
                                              end else begin
                                                if (6'h39 == _T_223) begin
                                                  mem_57 <= _GEN_14;
                                                end else begin
                                                  if (6'h39 == _T_218) begin
                                                    mem_57 <= _GEN_13;
                                                  end else begin
                                                    if (6'h39 == _T_213) begin
                                                      mem_57 <= _GEN_12;
                                                    end else begin
                                                      if (6'h39 == _T_208) begin
                                                        mem_57 <= _GEN_11;
                                                      end else begin
                                                        if (6'h39 == _T_203) begin
                                                          mem_57 <= _GEN_10;
                                                        end else begin
                                                          if (6'h39 == _T_198) begin
                                                            mem_57 <= _GEN_9;
                                                          end else begin
                                                            if (6'h39 == _T_193) begin
                                                              mem_57 <= _GEN_8;
                                                            end else begin
                                                              if (6'h39 == _T_188) begin
                                                                mem_57 <= _GEN_7;
                                                              end else begin
                                                                if (6'h39 == _T_183) begin
                                                                  mem_57 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h39 == _T_178) begin
                                                                    mem_57 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h39 == _T_173) begin
                                                                      mem_57 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h39 == _T_168) begin
                                                                        mem_57 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h39 == _T_163) begin
                                                                          mem_57 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h39 == _T_158) begin
                                                                            mem_57 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h39 == _T_153) begin
                                                                              mem_57 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h39 == _T_308) begin
              mem_57 <= _GEN_31;
            end else begin
              if (6'h39 == _T_303) begin
                mem_57 <= _GEN_30;
              end else begin
                if (6'h39 == _T_298) begin
                  mem_57 <= _GEN_29;
                end else begin
                  if (6'h39 == _T_293) begin
                    mem_57 <= _GEN_28;
                  end else begin
                    if (6'h39 == _T_288) begin
                      mem_57 <= _GEN_27;
                    end else begin
                      if (6'h39 == _T_283) begin
                        mem_57 <= _GEN_26;
                      end else begin
                        if (6'h39 == _T_278) begin
                          mem_57 <= _GEN_25;
                        end else begin
                          if (6'h39 == _T_273) begin
                            mem_57 <= _GEN_24;
                          end else begin
                            if (6'h39 == _T_268) begin
                              mem_57 <= _GEN_23;
                            end else begin
                              if (6'h39 == _T_263) begin
                                mem_57 <= _GEN_22;
                              end else begin
                                if (6'h39 == _T_258) begin
                                  mem_57 <= _GEN_21;
                                end else begin
                                  if (6'h39 == _T_253) begin
                                    mem_57 <= _GEN_20;
                                  end else begin
                                    if (6'h39 == _T_248) begin
                                      mem_57 <= _GEN_19;
                                    end else begin
                                      if (6'h39 == _T_243) begin
                                        mem_57 <= _GEN_18;
                                      end else begin
                                        if (6'h39 == _T_238) begin
                                          mem_57 <= _GEN_17;
                                        end else begin
                                          if (6'h39 == _T_233) begin
                                            mem_57 <= _GEN_16;
                                          end else begin
                                            if (6'h39 == _T_228) begin
                                              mem_57 <= _GEN_15;
                                            end else begin
                                              if (6'h39 == _T_223) begin
                                                mem_57 <= _GEN_14;
                                              end else begin
                                                if (6'h39 == _T_218) begin
                                                  mem_57 <= _GEN_13;
                                                end else begin
                                                  if (6'h39 == _T_213) begin
                                                    mem_57 <= _GEN_12;
                                                  end else begin
                                                    if (6'h39 == _T_208) begin
                                                      mem_57 <= _GEN_11;
                                                    end else begin
                                                      if (6'h39 == _T_203) begin
                                                        mem_57 <= _GEN_10;
                                                      end else begin
                                                        if (6'h39 == _T_198) begin
                                                          mem_57 <= _GEN_9;
                                                        end else begin
                                                          if (6'h39 == _T_193) begin
                                                            mem_57 <= _GEN_8;
                                                          end else begin
                                                            if (6'h39 == _T_188) begin
                                                              mem_57 <= _GEN_7;
                                                            end else begin
                                                              if (6'h39 == _T_183) begin
                                                                mem_57 <= _GEN_6;
                                                              end else begin
                                                                if (6'h39 == _T_178) begin
                                                                  mem_57 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h39 == _T_173) begin
                                                                    mem_57 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h39 == _T_168) begin
                                                                      mem_57 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h39 == _T_163) begin
                                                                        mem_57 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h39 == _T_158) begin
                                                                          mem_57 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h39 == _T_153) begin
                                                                            mem_57 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h39 == _T_308) begin
            mem_57 <= _GEN_31;
          end else begin
            if (6'h39 == _T_303) begin
              mem_57 <= _GEN_30;
            end else begin
              if (6'h39 == _T_298) begin
                mem_57 <= _GEN_29;
              end else begin
                if (6'h39 == _T_293) begin
                  mem_57 <= _GEN_28;
                end else begin
                  if (6'h39 == _T_288) begin
                    mem_57 <= _GEN_27;
                  end else begin
                    if (6'h39 == _T_283) begin
                      mem_57 <= _GEN_26;
                    end else begin
                      if (6'h39 == _T_278) begin
                        mem_57 <= _GEN_25;
                      end else begin
                        if (6'h39 == _T_273) begin
                          mem_57 <= _GEN_24;
                        end else begin
                          if (6'h39 == _T_268) begin
                            mem_57 <= _GEN_23;
                          end else begin
                            if (6'h39 == _T_263) begin
                              mem_57 <= _GEN_22;
                            end else begin
                              if (6'h39 == _T_258) begin
                                mem_57 <= _GEN_21;
                              end else begin
                                if (6'h39 == _T_253) begin
                                  mem_57 <= _GEN_20;
                                end else begin
                                  if (6'h39 == _T_248) begin
                                    mem_57 <= _GEN_19;
                                  end else begin
                                    if (6'h39 == _T_243) begin
                                      mem_57 <= _GEN_18;
                                    end else begin
                                      if (6'h39 == _T_238) begin
                                        mem_57 <= _GEN_17;
                                      end else begin
                                        if (6'h39 == _T_233) begin
                                          mem_57 <= _GEN_16;
                                        end else begin
                                          if (6'h39 == _T_228) begin
                                            mem_57 <= _GEN_15;
                                          end else begin
                                            if (6'h39 == _T_223) begin
                                              mem_57 <= _GEN_14;
                                            end else begin
                                              if (6'h39 == _T_218) begin
                                                mem_57 <= _GEN_13;
                                              end else begin
                                                if (6'h39 == _T_213) begin
                                                  mem_57 <= _GEN_12;
                                                end else begin
                                                  if (6'h39 == _T_208) begin
                                                    mem_57 <= _GEN_11;
                                                  end else begin
                                                    if (6'h39 == _T_203) begin
                                                      mem_57 <= _GEN_10;
                                                    end else begin
                                                      if (6'h39 == _T_198) begin
                                                        mem_57 <= _GEN_9;
                                                      end else begin
                                                        if (6'h39 == _T_193) begin
                                                          mem_57 <= _GEN_8;
                                                        end else begin
                                                          if (6'h39 == _T_188) begin
                                                            mem_57 <= _GEN_7;
                                                          end else begin
                                                            if (6'h39 == _T_183) begin
                                                              mem_57 <= _GEN_6;
                                                            end else begin
                                                              if (6'h39 == _T_178) begin
                                                                mem_57 <= _GEN_5;
                                                              end else begin
                                                                if (6'h39 == _T_173) begin
                                                                  mem_57 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h39 == _T_168) begin
                                                                    mem_57 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h39 == _T_163) begin
                                                                      mem_57 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h39 == _T_158) begin
                                                                        mem_57 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h39 == _T_153) begin
                                                                          mem_57 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h39 == _T_308) begin
          mem_57 <= _GEN_31;
        end else begin
          if (6'h39 == _T_303) begin
            mem_57 <= _GEN_30;
          end else begin
            if (6'h39 == _T_298) begin
              mem_57 <= _GEN_29;
            end else begin
              if (6'h39 == _T_293) begin
                mem_57 <= _GEN_28;
              end else begin
                if (6'h39 == _T_288) begin
                  mem_57 <= _GEN_27;
                end else begin
                  if (6'h39 == _T_283) begin
                    mem_57 <= _GEN_26;
                  end else begin
                    if (6'h39 == _T_278) begin
                      mem_57 <= _GEN_25;
                    end else begin
                      if (6'h39 == _T_273) begin
                        mem_57 <= _GEN_24;
                      end else begin
                        if (6'h39 == _T_268) begin
                          mem_57 <= _GEN_23;
                        end else begin
                          if (6'h39 == _T_263) begin
                            mem_57 <= _GEN_22;
                          end else begin
                            if (6'h39 == _T_258) begin
                              mem_57 <= _GEN_21;
                            end else begin
                              if (6'h39 == _T_253) begin
                                mem_57 <= _GEN_20;
                              end else begin
                                if (6'h39 == _T_248) begin
                                  mem_57 <= _GEN_19;
                                end else begin
                                  if (6'h39 == _T_243) begin
                                    mem_57 <= _GEN_18;
                                  end else begin
                                    if (6'h39 == _T_238) begin
                                      mem_57 <= _GEN_17;
                                    end else begin
                                      if (6'h39 == _T_233) begin
                                        mem_57 <= _GEN_16;
                                      end else begin
                                        if (6'h39 == _T_228) begin
                                          mem_57 <= _GEN_15;
                                        end else begin
                                          if (6'h39 == _T_223) begin
                                            mem_57 <= _GEN_14;
                                          end else begin
                                            if (6'h39 == _T_218) begin
                                              mem_57 <= _GEN_13;
                                            end else begin
                                              if (6'h39 == _T_213) begin
                                                mem_57 <= _GEN_12;
                                              end else begin
                                                if (6'h39 == _T_208) begin
                                                  mem_57 <= _GEN_11;
                                                end else begin
                                                  if (6'h39 == _T_203) begin
                                                    mem_57 <= _GEN_10;
                                                  end else begin
                                                    if (6'h39 == _T_198) begin
                                                      mem_57 <= _GEN_9;
                                                    end else begin
                                                      if (6'h39 == _T_193) begin
                                                        mem_57 <= _GEN_8;
                                                      end else begin
                                                        if (6'h39 == _T_188) begin
                                                          mem_57 <= _GEN_7;
                                                        end else begin
                                                          if (6'h39 == _T_183) begin
                                                            mem_57 <= _GEN_6;
                                                          end else begin
                                                            if (6'h39 == _T_178) begin
                                                              mem_57 <= _GEN_5;
                                                            end else begin
                                                              if (6'h39 == _T_173) begin
                                                                mem_57 <= _GEN_4;
                                                              end else begin
                                                                if (6'h39 == _T_168) begin
                                                                  mem_57 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h39 == _T_163) begin
                                                                    mem_57 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h39 == _T_158) begin
                                                                      mem_57 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h39 == _T_153) begin
                                                                        mem_57 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h3a == wPos) begin
            mem_58 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h3a == _T_308) begin
                mem_58 <= _GEN_31;
              end else begin
                if (6'h3a == _T_303) begin
                  mem_58 <= _GEN_30;
                end else begin
                  if (6'h3a == _T_298) begin
                    mem_58 <= _GEN_29;
                  end else begin
                    if (6'h3a == _T_293) begin
                      mem_58 <= _GEN_28;
                    end else begin
                      if (6'h3a == _T_288) begin
                        mem_58 <= _GEN_27;
                      end else begin
                        if (6'h3a == _T_283) begin
                          mem_58 <= _GEN_26;
                        end else begin
                          if (6'h3a == _T_278) begin
                            mem_58 <= _GEN_25;
                          end else begin
                            if (6'h3a == _T_273) begin
                              mem_58 <= _GEN_24;
                            end else begin
                              if (6'h3a == _T_268) begin
                                mem_58 <= _GEN_23;
                              end else begin
                                if (6'h3a == _T_263) begin
                                  mem_58 <= _GEN_22;
                                end else begin
                                  if (6'h3a == _T_258) begin
                                    mem_58 <= _GEN_21;
                                  end else begin
                                    if (6'h3a == _T_253) begin
                                      mem_58 <= _GEN_20;
                                    end else begin
                                      if (6'h3a == _T_248) begin
                                        mem_58 <= _GEN_19;
                                      end else begin
                                        if (6'h3a == _T_243) begin
                                          mem_58 <= _GEN_18;
                                        end else begin
                                          if (6'h3a == _T_238) begin
                                            mem_58 <= _GEN_17;
                                          end else begin
                                            if (6'h3a == _T_233) begin
                                              mem_58 <= _GEN_16;
                                            end else begin
                                              if (6'h3a == _T_228) begin
                                                mem_58 <= _GEN_15;
                                              end else begin
                                                if (6'h3a == _T_223) begin
                                                  mem_58 <= _GEN_14;
                                                end else begin
                                                  if (6'h3a == _T_218) begin
                                                    mem_58 <= _GEN_13;
                                                  end else begin
                                                    if (6'h3a == _T_213) begin
                                                      mem_58 <= _GEN_12;
                                                    end else begin
                                                      if (6'h3a == _T_208) begin
                                                        mem_58 <= _GEN_11;
                                                      end else begin
                                                        if (6'h3a == _T_203) begin
                                                          mem_58 <= _GEN_10;
                                                        end else begin
                                                          if (6'h3a == _T_198) begin
                                                            mem_58 <= _GEN_9;
                                                          end else begin
                                                            if (6'h3a == _T_193) begin
                                                              mem_58 <= _GEN_8;
                                                            end else begin
                                                              if (6'h3a == _T_188) begin
                                                                mem_58 <= _GEN_7;
                                                              end else begin
                                                                if (6'h3a == _T_183) begin
                                                                  mem_58 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h3a == _T_178) begin
                                                                    mem_58 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h3a == _T_173) begin
                                                                      mem_58 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h3a == _T_168) begin
                                                                        mem_58 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h3a == _T_163) begin
                                                                          mem_58 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h3a == _T_158) begin
                                                                            mem_58 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h3a == _T_153) begin
                                                                              mem_58 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h3a == _T_308) begin
              mem_58 <= _GEN_31;
            end else begin
              if (6'h3a == _T_303) begin
                mem_58 <= _GEN_30;
              end else begin
                if (6'h3a == _T_298) begin
                  mem_58 <= _GEN_29;
                end else begin
                  if (6'h3a == _T_293) begin
                    mem_58 <= _GEN_28;
                  end else begin
                    if (6'h3a == _T_288) begin
                      mem_58 <= _GEN_27;
                    end else begin
                      if (6'h3a == _T_283) begin
                        mem_58 <= _GEN_26;
                      end else begin
                        if (6'h3a == _T_278) begin
                          mem_58 <= _GEN_25;
                        end else begin
                          if (6'h3a == _T_273) begin
                            mem_58 <= _GEN_24;
                          end else begin
                            if (6'h3a == _T_268) begin
                              mem_58 <= _GEN_23;
                            end else begin
                              if (6'h3a == _T_263) begin
                                mem_58 <= _GEN_22;
                              end else begin
                                if (6'h3a == _T_258) begin
                                  mem_58 <= _GEN_21;
                                end else begin
                                  if (6'h3a == _T_253) begin
                                    mem_58 <= _GEN_20;
                                  end else begin
                                    if (6'h3a == _T_248) begin
                                      mem_58 <= _GEN_19;
                                    end else begin
                                      if (6'h3a == _T_243) begin
                                        mem_58 <= _GEN_18;
                                      end else begin
                                        if (6'h3a == _T_238) begin
                                          mem_58 <= _GEN_17;
                                        end else begin
                                          if (6'h3a == _T_233) begin
                                            mem_58 <= _GEN_16;
                                          end else begin
                                            if (6'h3a == _T_228) begin
                                              mem_58 <= _GEN_15;
                                            end else begin
                                              if (6'h3a == _T_223) begin
                                                mem_58 <= _GEN_14;
                                              end else begin
                                                if (6'h3a == _T_218) begin
                                                  mem_58 <= _GEN_13;
                                                end else begin
                                                  if (6'h3a == _T_213) begin
                                                    mem_58 <= _GEN_12;
                                                  end else begin
                                                    if (6'h3a == _T_208) begin
                                                      mem_58 <= _GEN_11;
                                                    end else begin
                                                      if (6'h3a == _T_203) begin
                                                        mem_58 <= _GEN_10;
                                                      end else begin
                                                        if (6'h3a == _T_198) begin
                                                          mem_58 <= _GEN_9;
                                                        end else begin
                                                          if (6'h3a == _T_193) begin
                                                            mem_58 <= _GEN_8;
                                                          end else begin
                                                            if (6'h3a == _T_188) begin
                                                              mem_58 <= _GEN_7;
                                                            end else begin
                                                              if (6'h3a == _T_183) begin
                                                                mem_58 <= _GEN_6;
                                                              end else begin
                                                                if (6'h3a == _T_178) begin
                                                                  mem_58 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h3a == _T_173) begin
                                                                    mem_58 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h3a == _T_168) begin
                                                                      mem_58 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h3a == _T_163) begin
                                                                        mem_58 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h3a == _T_158) begin
                                                                          mem_58 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h3a == _T_153) begin
                                                                            mem_58 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h3a == _T_308) begin
            mem_58 <= _GEN_31;
          end else begin
            if (6'h3a == _T_303) begin
              mem_58 <= _GEN_30;
            end else begin
              if (6'h3a == _T_298) begin
                mem_58 <= _GEN_29;
              end else begin
                if (6'h3a == _T_293) begin
                  mem_58 <= _GEN_28;
                end else begin
                  if (6'h3a == _T_288) begin
                    mem_58 <= _GEN_27;
                  end else begin
                    if (6'h3a == _T_283) begin
                      mem_58 <= _GEN_26;
                    end else begin
                      if (6'h3a == _T_278) begin
                        mem_58 <= _GEN_25;
                      end else begin
                        if (6'h3a == _T_273) begin
                          mem_58 <= _GEN_24;
                        end else begin
                          if (6'h3a == _T_268) begin
                            mem_58 <= _GEN_23;
                          end else begin
                            if (6'h3a == _T_263) begin
                              mem_58 <= _GEN_22;
                            end else begin
                              if (6'h3a == _T_258) begin
                                mem_58 <= _GEN_21;
                              end else begin
                                if (6'h3a == _T_253) begin
                                  mem_58 <= _GEN_20;
                                end else begin
                                  if (6'h3a == _T_248) begin
                                    mem_58 <= _GEN_19;
                                  end else begin
                                    if (6'h3a == _T_243) begin
                                      mem_58 <= _GEN_18;
                                    end else begin
                                      if (6'h3a == _T_238) begin
                                        mem_58 <= _GEN_17;
                                      end else begin
                                        if (6'h3a == _T_233) begin
                                          mem_58 <= _GEN_16;
                                        end else begin
                                          if (6'h3a == _T_228) begin
                                            mem_58 <= _GEN_15;
                                          end else begin
                                            if (6'h3a == _T_223) begin
                                              mem_58 <= _GEN_14;
                                            end else begin
                                              if (6'h3a == _T_218) begin
                                                mem_58 <= _GEN_13;
                                              end else begin
                                                if (6'h3a == _T_213) begin
                                                  mem_58 <= _GEN_12;
                                                end else begin
                                                  if (6'h3a == _T_208) begin
                                                    mem_58 <= _GEN_11;
                                                  end else begin
                                                    if (6'h3a == _T_203) begin
                                                      mem_58 <= _GEN_10;
                                                    end else begin
                                                      if (6'h3a == _T_198) begin
                                                        mem_58 <= _GEN_9;
                                                      end else begin
                                                        if (6'h3a == _T_193) begin
                                                          mem_58 <= _GEN_8;
                                                        end else begin
                                                          if (6'h3a == _T_188) begin
                                                            mem_58 <= _GEN_7;
                                                          end else begin
                                                            if (6'h3a == _T_183) begin
                                                              mem_58 <= _GEN_6;
                                                            end else begin
                                                              if (6'h3a == _T_178) begin
                                                                mem_58 <= _GEN_5;
                                                              end else begin
                                                                if (6'h3a == _T_173) begin
                                                                  mem_58 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h3a == _T_168) begin
                                                                    mem_58 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h3a == _T_163) begin
                                                                      mem_58 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h3a == _T_158) begin
                                                                        mem_58 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h3a == _T_153) begin
                                                                          mem_58 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h3a == _T_308) begin
          mem_58 <= _GEN_31;
        end else begin
          if (6'h3a == _T_303) begin
            mem_58 <= _GEN_30;
          end else begin
            if (6'h3a == _T_298) begin
              mem_58 <= _GEN_29;
            end else begin
              if (6'h3a == _T_293) begin
                mem_58 <= _GEN_28;
              end else begin
                if (6'h3a == _T_288) begin
                  mem_58 <= _GEN_27;
                end else begin
                  if (6'h3a == _T_283) begin
                    mem_58 <= _GEN_26;
                  end else begin
                    if (6'h3a == _T_278) begin
                      mem_58 <= _GEN_25;
                    end else begin
                      if (6'h3a == _T_273) begin
                        mem_58 <= _GEN_24;
                      end else begin
                        if (6'h3a == _T_268) begin
                          mem_58 <= _GEN_23;
                        end else begin
                          if (6'h3a == _T_263) begin
                            mem_58 <= _GEN_22;
                          end else begin
                            if (6'h3a == _T_258) begin
                              mem_58 <= _GEN_21;
                            end else begin
                              if (6'h3a == _T_253) begin
                                mem_58 <= _GEN_20;
                              end else begin
                                if (6'h3a == _T_248) begin
                                  mem_58 <= _GEN_19;
                                end else begin
                                  if (6'h3a == _T_243) begin
                                    mem_58 <= _GEN_18;
                                  end else begin
                                    if (6'h3a == _T_238) begin
                                      mem_58 <= _GEN_17;
                                    end else begin
                                      if (6'h3a == _T_233) begin
                                        mem_58 <= _GEN_16;
                                      end else begin
                                        if (6'h3a == _T_228) begin
                                          mem_58 <= _GEN_15;
                                        end else begin
                                          if (6'h3a == _T_223) begin
                                            mem_58 <= _GEN_14;
                                          end else begin
                                            if (6'h3a == _T_218) begin
                                              mem_58 <= _GEN_13;
                                            end else begin
                                              if (6'h3a == _T_213) begin
                                                mem_58 <= _GEN_12;
                                              end else begin
                                                if (6'h3a == _T_208) begin
                                                  mem_58 <= _GEN_11;
                                                end else begin
                                                  if (6'h3a == _T_203) begin
                                                    mem_58 <= _GEN_10;
                                                  end else begin
                                                    if (6'h3a == _T_198) begin
                                                      mem_58 <= _GEN_9;
                                                    end else begin
                                                      if (6'h3a == _T_193) begin
                                                        mem_58 <= _GEN_8;
                                                      end else begin
                                                        if (6'h3a == _T_188) begin
                                                          mem_58 <= _GEN_7;
                                                        end else begin
                                                          if (6'h3a == _T_183) begin
                                                            mem_58 <= _GEN_6;
                                                          end else begin
                                                            if (6'h3a == _T_178) begin
                                                              mem_58 <= _GEN_5;
                                                            end else begin
                                                              if (6'h3a == _T_173) begin
                                                                mem_58 <= _GEN_4;
                                                              end else begin
                                                                if (6'h3a == _T_168) begin
                                                                  mem_58 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h3a == _T_163) begin
                                                                    mem_58 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h3a == _T_158) begin
                                                                      mem_58 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h3a == _T_153) begin
                                                                        mem_58 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h3b == wPos) begin
            mem_59 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h3b == _T_308) begin
                mem_59 <= _GEN_31;
              end else begin
                if (6'h3b == _T_303) begin
                  mem_59 <= _GEN_30;
                end else begin
                  if (6'h3b == _T_298) begin
                    mem_59 <= _GEN_29;
                  end else begin
                    if (6'h3b == _T_293) begin
                      mem_59 <= _GEN_28;
                    end else begin
                      if (6'h3b == _T_288) begin
                        mem_59 <= _GEN_27;
                      end else begin
                        if (6'h3b == _T_283) begin
                          mem_59 <= _GEN_26;
                        end else begin
                          if (6'h3b == _T_278) begin
                            mem_59 <= _GEN_25;
                          end else begin
                            if (6'h3b == _T_273) begin
                              mem_59 <= _GEN_24;
                            end else begin
                              if (6'h3b == _T_268) begin
                                mem_59 <= _GEN_23;
                              end else begin
                                if (6'h3b == _T_263) begin
                                  mem_59 <= _GEN_22;
                                end else begin
                                  if (6'h3b == _T_258) begin
                                    mem_59 <= _GEN_21;
                                  end else begin
                                    if (6'h3b == _T_253) begin
                                      mem_59 <= _GEN_20;
                                    end else begin
                                      if (6'h3b == _T_248) begin
                                        mem_59 <= _GEN_19;
                                      end else begin
                                        if (6'h3b == _T_243) begin
                                          mem_59 <= _GEN_18;
                                        end else begin
                                          if (6'h3b == _T_238) begin
                                            mem_59 <= _GEN_17;
                                          end else begin
                                            if (6'h3b == _T_233) begin
                                              mem_59 <= _GEN_16;
                                            end else begin
                                              if (6'h3b == _T_228) begin
                                                mem_59 <= _GEN_15;
                                              end else begin
                                                if (6'h3b == _T_223) begin
                                                  mem_59 <= _GEN_14;
                                                end else begin
                                                  if (6'h3b == _T_218) begin
                                                    mem_59 <= _GEN_13;
                                                  end else begin
                                                    if (6'h3b == _T_213) begin
                                                      mem_59 <= _GEN_12;
                                                    end else begin
                                                      if (6'h3b == _T_208) begin
                                                        mem_59 <= _GEN_11;
                                                      end else begin
                                                        if (6'h3b == _T_203) begin
                                                          mem_59 <= _GEN_10;
                                                        end else begin
                                                          if (6'h3b == _T_198) begin
                                                            mem_59 <= _GEN_9;
                                                          end else begin
                                                            if (6'h3b == _T_193) begin
                                                              mem_59 <= _GEN_8;
                                                            end else begin
                                                              if (6'h3b == _T_188) begin
                                                                mem_59 <= _GEN_7;
                                                              end else begin
                                                                if (6'h3b == _T_183) begin
                                                                  mem_59 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h3b == _T_178) begin
                                                                    mem_59 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h3b == _T_173) begin
                                                                      mem_59 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h3b == _T_168) begin
                                                                        mem_59 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h3b == _T_163) begin
                                                                          mem_59 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h3b == _T_158) begin
                                                                            mem_59 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h3b == _T_153) begin
                                                                              mem_59 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h3b == _T_308) begin
              mem_59 <= _GEN_31;
            end else begin
              if (6'h3b == _T_303) begin
                mem_59 <= _GEN_30;
              end else begin
                if (6'h3b == _T_298) begin
                  mem_59 <= _GEN_29;
                end else begin
                  if (6'h3b == _T_293) begin
                    mem_59 <= _GEN_28;
                  end else begin
                    if (6'h3b == _T_288) begin
                      mem_59 <= _GEN_27;
                    end else begin
                      if (6'h3b == _T_283) begin
                        mem_59 <= _GEN_26;
                      end else begin
                        if (6'h3b == _T_278) begin
                          mem_59 <= _GEN_25;
                        end else begin
                          if (6'h3b == _T_273) begin
                            mem_59 <= _GEN_24;
                          end else begin
                            if (6'h3b == _T_268) begin
                              mem_59 <= _GEN_23;
                            end else begin
                              if (6'h3b == _T_263) begin
                                mem_59 <= _GEN_22;
                              end else begin
                                if (6'h3b == _T_258) begin
                                  mem_59 <= _GEN_21;
                                end else begin
                                  if (6'h3b == _T_253) begin
                                    mem_59 <= _GEN_20;
                                  end else begin
                                    if (6'h3b == _T_248) begin
                                      mem_59 <= _GEN_19;
                                    end else begin
                                      if (6'h3b == _T_243) begin
                                        mem_59 <= _GEN_18;
                                      end else begin
                                        if (6'h3b == _T_238) begin
                                          mem_59 <= _GEN_17;
                                        end else begin
                                          if (6'h3b == _T_233) begin
                                            mem_59 <= _GEN_16;
                                          end else begin
                                            if (6'h3b == _T_228) begin
                                              mem_59 <= _GEN_15;
                                            end else begin
                                              if (6'h3b == _T_223) begin
                                                mem_59 <= _GEN_14;
                                              end else begin
                                                if (6'h3b == _T_218) begin
                                                  mem_59 <= _GEN_13;
                                                end else begin
                                                  if (6'h3b == _T_213) begin
                                                    mem_59 <= _GEN_12;
                                                  end else begin
                                                    if (6'h3b == _T_208) begin
                                                      mem_59 <= _GEN_11;
                                                    end else begin
                                                      if (6'h3b == _T_203) begin
                                                        mem_59 <= _GEN_10;
                                                      end else begin
                                                        if (6'h3b == _T_198) begin
                                                          mem_59 <= _GEN_9;
                                                        end else begin
                                                          if (6'h3b == _T_193) begin
                                                            mem_59 <= _GEN_8;
                                                          end else begin
                                                            if (6'h3b == _T_188) begin
                                                              mem_59 <= _GEN_7;
                                                            end else begin
                                                              if (6'h3b == _T_183) begin
                                                                mem_59 <= _GEN_6;
                                                              end else begin
                                                                if (6'h3b == _T_178) begin
                                                                  mem_59 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h3b == _T_173) begin
                                                                    mem_59 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h3b == _T_168) begin
                                                                      mem_59 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h3b == _T_163) begin
                                                                        mem_59 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h3b == _T_158) begin
                                                                          mem_59 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h3b == _T_153) begin
                                                                            mem_59 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h3b == _T_308) begin
            mem_59 <= _GEN_31;
          end else begin
            if (6'h3b == _T_303) begin
              mem_59 <= _GEN_30;
            end else begin
              if (6'h3b == _T_298) begin
                mem_59 <= _GEN_29;
              end else begin
                if (6'h3b == _T_293) begin
                  mem_59 <= _GEN_28;
                end else begin
                  if (6'h3b == _T_288) begin
                    mem_59 <= _GEN_27;
                  end else begin
                    if (6'h3b == _T_283) begin
                      mem_59 <= _GEN_26;
                    end else begin
                      if (6'h3b == _T_278) begin
                        mem_59 <= _GEN_25;
                      end else begin
                        if (6'h3b == _T_273) begin
                          mem_59 <= _GEN_24;
                        end else begin
                          if (6'h3b == _T_268) begin
                            mem_59 <= _GEN_23;
                          end else begin
                            if (6'h3b == _T_263) begin
                              mem_59 <= _GEN_22;
                            end else begin
                              if (6'h3b == _T_258) begin
                                mem_59 <= _GEN_21;
                              end else begin
                                if (6'h3b == _T_253) begin
                                  mem_59 <= _GEN_20;
                                end else begin
                                  if (6'h3b == _T_248) begin
                                    mem_59 <= _GEN_19;
                                  end else begin
                                    if (6'h3b == _T_243) begin
                                      mem_59 <= _GEN_18;
                                    end else begin
                                      if (6'h3b == _T_238) begin
                                        mem_59 <= _GEN_17;
                                      end else begin
                                        if (6'h3b == _T_233) begin
                                          mem_59 <= _GEN_16;
                                        end else begin
                                          if (6'h3b == _T_228) begin
                                            mem_59 <= _GEN_15;
                                          end else begin
                                            if (6'h3b == _T_223) begin
                                              mem_59 <= _GEN_14;
                                            end else begin
                                              if (6'h3b == _T_218) begin
                                                mem_59 <= _GEN_13;
                                              end else begin
                                                if (6'h3b == _T_213) begin
                                                  mem_59 <= _GEN_12;
                                                end else begin
                                                  if (6'h3b == _T_208) begin
                                                    mem_59 <= _GEN_11;
                                                  end else begin
                                                    if (6'h3b == _T_203) begin
                                                      mem_59 <= _GEN_10;
                                                    end else begin
                                                      if (6'h3b == _T_198) begin
                                                        mem_59 <= _GEN_9;
                                                      end else begin
                                                        if (6'h3b == _T_193) begin
                                                          mem_59 <= _GEN_8;
                                                        end else begin
                                                          if (6'h3b == _T_188) begin
                                                            mem_59 <= _GEN_7;
                                                          end else begin
                                                            if (6'h3b == _T_183) begin
                                                              mem_59 <= _GEN_6;
                                                            end else begin
                                                              if (6'h3b == _T_178) begin
                                                                mem_59 <= _GEN_5;
                                                              end else begin
                                                                if (6'h3b == _T_173) begin
                                                                  mem_59 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h3b == _T_168) begin
                                                                    mem_59 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h3b == _T_163) begin
                                                                      mem_59 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h3b == _T_158) begin
                                                                        mem_59 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h3b == _T_153) begin
                                                                          mem_59 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h3b == _T_308) begin
          mem_59 <= _GEN_31;
        end else begin
          if (6'h3b == _T_303) begin
            mem_59 <= _GEN_30;
          end else begin
            if (6'h3b == _T_298) begin
              mem_59 <= _GEN_29;
            end else begin
              if (6'h3b == _T_293) begin
                mem_59 <= _GEN_28;
              end else begin
                if (6'h3b == _T_288) begin
                  mem_59 <= _GEN_27;
                end else begin
                  if (6'h3b == _T_283) begin
                    mem_59 <= _GEN_26;
                  end else begin
                    if (6'h3b == _T_278) begin
                      mem_59 <= _GEN_25;
                    end else begin
                      if (6'h3b == _T_273) begin
                        mem_59 <= _GEN_24;
                      end else begin
                        if (6'h3b == _T_268) begin
                          mem_59 <= _GEN_23;
                        end else begin
                          if (6'h3b == _T_263) begin
                            mem_59 <= _GEN_22;
                          end else begin
                            if (6'h3b == _T_258) begin
                              mem_59 <= _GEN_21;
                            end else begin
                              if (6'h3b == _T_253) begin
                                mem_59 <= _GEN_20;
                              end else begin
                                if (6'h3b == _T_248) begin
                                  mem_59 <= _GEN_19;
                                end else begin
                                  if (6'h3b == _T_243) begin
                                    mem_59 <= _GEN_18;
                                  end else begin
                                    if (6'h3b == _T_238) begin
                                      mem_59 <= _GEN_17;
                                    end else begin
                                      if (6'h3b == _T_233) begin
                                        mem_59 <= _GEN_16;
                                      end else begin
                                        if (6'h3b == _T_228) begin
                                          mem_59 <= _GEN_15;
                                        end else begin
                                          if (6'h3b == _T_223) begin
                                            mem_59 <= _GEN_14;
                                          end else begin
                                            if (6'h3b == _T_218) begin
                                              mem_59 <= _GEN_13;
                                            end else begin
                                              if (6'h3b == _T_213) begin
                                                mem_59 <= _GEN_12;
                                              end else begin
                                                if (6'h3b == _T_208) begin
                                                  mem_59 <= _GEN_11;
                                                end else begin
                                                  if (6'h3b == _T_203) begin
                                                    mem_59 <= _GEN_10;
                                                  end else begin
                                                    if (6'h3b == _T_198) begin
                                                      mem_59 <= _GEN_9;
                                                    end else begin
                                                      if (6'h3b == _T_193) begin
                                                        mem_59 <= _GEN_8;
                                                      end else begin
                                                        if (6'h3b == _T_188) begin
                                                          mem_59 <= _GEN_7;
                                                        end else begin
                                                          if (6'h3b == _T_183) begin
                                                            mem_59 <= _GEN_6;
                                                          end else begin
                                                            if (6'h3b == _T_178) begin
                                                              mem_59 <= _GEN_5;
                                                            end else begin
                                                              if (6'h3b == _T_173) begin
                                                                mem_59 <= _GEN_4;
                                                              end else begin
                                                                if (6'h3b == _T_168) begin
                                                                  mem_59 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h3b == _T_163) begin
                                                                    mem_59 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h3b == _T_158) begin
                                                                      mem_59 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h3b == _T_153) begin
                                                                        mem_59 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h3c == wPos) begin
            mem_60 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h3c == _T_308) begin
                mem_60 <= _GEN_31;
              end else begin
                if (6'h3c == _T_303) begin
                  mem_60 <= _GEN_30;
                end else begin
                  if (6'h3c == _T_298) begin
                    mem_60 <= _GEN_29;
                  end else begin
                    if (6'h3c == _T_293) begin
                      mem_60 <= _GEN_28;
                    end else begin
                      if (6'h3c == _T_288) begin
                        mem_60 <= _GEN_27;
                      end else begin
                        if (6'h3c == _T_283) begin
                          mem_60 <= _GEN_26;
                        end else begin
                          if (6'h3c == _T_278) begin
                            mem_60 <= _GEN_25;
                          end else begin
                            if (6'h3c == _T_273) begin
                              mem_60 <= _GEN_24;
                            end else begin
                              if (6'h3c == _T_268) begin
                                mem_60 <= _GEN_23;
                              end else begin
                                if (6'h3c == _T_263) begin
                                  mem_60 <= _GEN_22;
                                end else begin
                                  if (6'h3c == _T_258) begin
                                    mem_60 <= _GEN_21;
                                  end else begin
                                    if (6'h3c == _T_253) begin
                                      mem_60 <= _GEN_20;
                                    end else begin
                                      if (6'h3c == _T_248) begin
                                        mem_60 <= _GEN_19;
                                      end else begin
                                        if (6'h3c == _T_243) begin
                                          mem_60 <= _GEN_18;
                                        end else begin
                                          if (6'h3c == _T_238) begin
                                            mem_60 <= _GEN_17;
                                          end else begin
                                            if (6'h3c == _T_233) begin
                                              mem_60 <= _GEN_16;
                                            end else begin
                                              if (6'h3c == _T_228) begin
                                                mem_60 <= _GEN_15;
                                              end else begin
                                                if (6'h3c == _T_223) begin
                                                  mem_60 <= _GEN_14;
                                                end else begin
                                                  if (6'h3c == _T_218) begin
                                                    mem_60 <= _GEN_13;
                                                  end else begin
                                                    if (6'h3c == _T_213) begin
                                                      mem_60 <= _GEN_12;
                                                    end else begin
                                                      if (6'h3c == _T_208) begin
                                                        mem_60 <= _GEN_11;
                                                      end else begin
                                                        if (6'h3c == _T_203) begin
                                                          mem_60 <= _GEN_10;
                                                        end else begin
                                                          if (6'h3c == _T_198) begin
                                                            mem_60 <= _GEN_9;
                                                          end else begin
                                                            if (6'h3c == _T_193) begin
                                                              mem_60 <= _GEN_8;
                                                            end else begin
                                                              if (6'h3c == _T_188) begin
                                                                mem_60 <= _GEN_7;
                                                              end else begin
                                                                if (6'h3c == _T_183) begin
                                                                  mem_60 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h3c == _T_178) begin
                                                                    mem_60 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h3c == _T_173) begin
                                                                      mem_60 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h3c == _T_168) begin
                                                                        mem_60 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h3c == _T_163) begin
                                                                          mem_60 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h3c == _T_158) begin
                                                                            mem_60 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h3c == _T_153) begin
                                                                              mem_60 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h3c == _T_308) begin
              mem_60 <= _GEN_31;
            end else begin
              if (6'h3c == _T_303) begin
                mem_60 <= _GEN_30;
              end else begin
                if (6'h3c == _T_298) begin
                  mem_60 <= _GEN_29;
                end else begin
                  if (6'h3c == _T_293) begin
                    mem_60 <= _GEN_28;
                  end else begin
                    if (6'h3c == _T_288) begin
                      mem_60 <= _GEN_27;
                    end else begin
                      if (6'h3c == _T_283) begin
                        mem_60 <= _GEN_26;
                      end else begin
                        if (6'h3c == _T_278) begin
                          mem_60 <= _GEN_25;
                        end else begin
                          if (6'h3c == _T_273) begin
                            mem_60 <= _GEN_24;
                          end else begin
                            if (6'h3c == _T_268) begin
                              mem_60 <= _GEN_23;
                            end else begin
                              if (6'h3c == _T_263) begin
                                mem_60 <= _GEN_22;
                              end else begin
                                if (6'h3c == _T_258) begin
                                  mem_60 <= _GEN_21;
                                end else begin
                                  if (6'h3c == _T_253) begin
                                    mem_60 <= _GEN_20;
                                  end else begin
                                    if (6'h3c == _T_248) begin
                                      mem_60 <= _GEN_19;
                                    end else begin
                                      if (6'h3c == _T_243) begin
                                        mem_60 <= _GEN_18;
                                      end else begin
                                        if (6'h3c == _T_238) begin
                                          mem_60 <= _GEN_17;
                                        end else begin
                                          if (6'h3c == _T_233) begin
                                            mem_60 <= _GEN_16;
                                          end else begin
                                            if (6'h3c == _T_228) begin
                                              mem_60 <= _GEN_15;
                                            end else begin
                                              if (6'h3c == _T_223) begin
                                                mem_60 <= _GEN_14;
                                              end else begin
                                                if (6'h3c == _T_218) begin
                                                  mem_60 <= _GEN_13;
                                                end else begin
                                                  if (6'h3c == _T_213) begin
                                                    mem_60 <= _GEN_12;
                                                  end else begin
                                                    if (6'h3c == _T_208) begin
                                                      mem_60 <= _GEN_11;
                                                    end else begin
                                                      if (6'h3c == _T_203) begin
                                                        mem_60 <= _GEN_10;
                                                      end else begin
                                                        if (6'h3c == _T_198) begin
                                                          mem_60 <= _GEN_9;
                                                        end else begin
                                                          if (6'h3c == _T_193) begin
                                                            mem_60 <= _GEN_8;
                                                          end else begin
                                                            if (6'h3c == _T_188) begin
                                                              mem_60 <= _GEN_7;
                                                            end else begin
                                                              if (6'h3c == _T_183) begin
                                                                mem_60 <= _GEN_6;
                                                              end else begin
                                                                if (6'h3c == _T_178) begin
                                                                  mem_60 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h3c == _T_173) begin
                                                                    mem_60 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h3c == _T_168) begin
                                                                      mem_60 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h3c == _T_163) begin
                                                                        mem_60 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h3c == _T_158) begin
                                                                          mem_60 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h3c == _T_153) begin
                                                                            mem_60 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h3c == _T_308) begin
            mem_60 <= _GEN_31;
          end else begin
            if (6'h3c == _T_303) begin
              mem_60 <= _GEN_30;
            end else begin
              if (6'h3c == _T_298) begin
                mem_60 <= _GEN_29;
              end else begin
                if (6'h3c == _T_293) begin
                  mem_60 <= _GEN_28;
                end else begin
                  if (6'h3c == _T_288) begin
                    mem_60 <= _GEN_27;
                  end else begin
                    if (6'h3c == _T_283) begin
                      mem_60 <= _GEN_26;
                    end else begin
                      if (6'h3c == _T_278) begin
                        mem_60 <= _GEN_25;
                      end else begin
                        if (6'h3c == _T_273) begin
                          mem_60 <= _GEN_24;
                        end else begin
                          if (6'h3c == _T_268) begin
                            mem_60 <= _GEN_23;
                          end else begin
                            if (6'h3c == _T_263) begin
                              mem_60 <= _GEN_22;
                            end else begin
                              if (6'h3c == _T_258) begin
                                mem_60 <= _GEN_21;
                              end else begin
                                if (6'h3c == _T_253) begin
                                  mem_60 <= _GEN_20;
                                end else begin
                                  if (6'h3c == _T_248) begin
                                    mem_60 <= _GEN_19;
                                  end else begin
                                    if (6'h3c == _T_243) begin
                                      mem_60 <= _GEN_18;
                                    end else begin
                                      if (6'h3c == _T_238) begin
                                        mem_60 <= _GEN_17;
                                      end else begin
                                        if (6'h3c == _T_233) begin
                                          mem_60 <= _GEN_16;
                                        end else begin
                                          if (6'h3c == _T_228) begin
                                            mem_60 <= _GEN_15;
                                          end else begin
                                            if (6'h3c == _T_223) begin
                                              mem_60 <= _GEN_14;
                                            end else begin
                                              if (6'h3c == _T_218) begin
                                                mem_60 <= _GEN_13;
                                              end else begin
                                                if (6'h3c == _T_213) begin
                                                  mem_60 <= _GEN_12;
                                                end else begin
                                                  if (6'h3c == _T_208) begin
                                                    mem_60 <= _GEN_11;
                                                  end else begin
                                                    if (6'h3c == _T_203) begin
                                                      mem_60 <= _GEN_10;
                                                    end else begin
                                                      if (6'h3c == _T_198) begin
                                                        mem_60 <= _GEN_9;
                                                      end else begin
                                                        if (6'h3c == _T_193) begin
                                                          mem_60 <= _GEN_8;
                                                        end else begin
                                                          if (6'h3c == _T_188) begin
                                                            mem_60 <= _GEN_7;
                                                          end else begin
                                                            if (6'h3c == _T_183) begin
                                                              mem_60 <= _GEN_6;
                                                            end else begin
                                                              if (6'h3c == _T_178) begin
                                                                mem_60 <= _GEN_5;
                                                              end else begin
                                                                if (6'h3c == _T_173) begin
                                                                  mem_60 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h3c == _T_168) begin
                                                                    mem_60 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h3c == _T_163) begin
                                                                      mem_60 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h3c == _T_158) begin
                                                                        mem_60 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h3c == _T_153) begin
                                                                          mem_60 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h3c == _T_308) begin
          mem_60 <= _GEN_31;
        end else begin
          if (6'h3c == _T_303) begin
            mem_60 <= _GEN_30;
          end else begin
            if (6'h3c == _T_298) begin
              mem_60 <= _GEN_29;
            end else begin
              if (6'h3c == _T_293) begin
                mem_60 <= _GEN_28;
              end else begin
                if (6'h3c == _T_288) begin
                  mem_60 <= _GEN_27;
                end else begin
                  if (6'h3c == _T_283) begin
                    mem_60 <= _GEN_26;
                  end else begin
                    if (6'h3c == _T_278) begin
                      mem_60 <= _GEN_25;
                    end else begin
                      if (6'h3c == _T_273) begin
                        mem_60 <= _GEN_24;
                      end else begin
                        if (6'h3c == _T_268) begin
                          mem_60 <= _GEN_23;
                        end else begin
                          if (6'h3c == _T_263) begin
                            mem_60 <= _GEN_22;
                          end else begin
                            if (6'h3c == _T_258) begin
                              mem_60 <= _GEN_21;
                            end else begin
                              if (6'h3c == _T_253) begin
                                mem_60 <= _GEN_20;
                              end else begin
                                if (6'h3c == _T_248) begin
                                  mem_60 <= _GEN_19;
                                end else begin
                                  if (6'h3c == _T_243) begin
                                    mem_60 <= _GEN_18;
                                  end else begin
                                    if (6'h3c == _T_238) begin
                                      mem_60 <= _GEN_17;
                                    end else begin
                                      if (6'h3c == _T_233) begin
                                        mem_60 <= _GEN_16;
                                      end else begin
                                        if (6'h3c == _T_228) begin
                                          mem_60 <= _GEN_15;
                                        end else begin
                                          if (6'h3c == _T_223) begin
                                            mem_60 <= _GEN_14;
                                          end else begin
                                            if (6'h3c == _T_218) begin
                                              mem_60 <= _GEN_13;
                                            end else begin
                                              if (6'h3c == _T_213) begin
                                                mem_60 <= _GEN_12;
                                              end else begin
                                                if (6'h3c == _T_208) begin
                                                  mem_60 <= _GEN_11;
                                                end else begin
                                                  if (6'h3c == _T_203) begin
                                                    mem_60 <= _GEN_10;
                                                  end else begin
                                                    if (6'h3c == _T_198) begin
                                                      mem_60 <= _GEN_9;
                                                    end else begin
                                                      if (6'h3c == _T_193) begin
                                                        mem_60 <= _GEN_8;
                                                      end else begin
                                                        if (6'h3c == _T_188) begin
                                                          mem_60 <= _GEN_7;
                                                        end else begin
                                                          if (6'h3c == _T_183) begin
                                                            mem_60 <= _GEN_6;
                                                          end else begin
                                                            if (6'h3c == _T_178) begin
                                                              mem_60 <= _GEN_5;
                                                            end else begin
                                                              if (6'h3c == _T_173) begin
                                                                mem_60 <= _GEN_4;
                                                              end else begin
                                                                if (6'h3c == _T_168) begin
                                                                  mem_60 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h3c == _T_163) begin
                                                                    mem_60 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h3c == _T_158) begin
                                                                      mem_60 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h3c == _T_153) begin
                                                                        mem_60 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h3d == wPos) begin
            mem_61 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h3d == _T_308) begin
                mem_61 <= _GEN_31;
              end else begin
                if (6'h3d == _T_303) begin
                  mem_61 <= _GEN_30;
                end else begin
                  if (6'h3d == _T_298) begin
                    mem_61 <= _GEN_29;
                  end else begin
                    if (6'h3d == _T_293) begin
                      mem_61 <= _GEN_28;
                    end else begin
                      if (6'h3d == _T_288) begin
                        mem_61 <= _GEN_27;
                      end else begin
                        if (6'h3d == _T_283) begin
                          mem_61 <= _GEN_26;
                        end else begin
                          if (6'h3d == _T_278) begin
                            mem_61 <= _GEN_25;
                          end else begin
                            if (6'h3d == _T_273) begin
                              mem_61 <= _GEN_24;
                            end else begin
                              if (6'h3d == _T_268) begin
                                mem_61 <= _GEN_23;
                              end else begin
                                if (6'h3d == _T_263) begin
                                  mem_61 <= _GEN_22;
                                end else begin
                                  if (6'h3d == _T_258) begin
                                    mem_61 <= _GEN_21;
                                  end else begin
                                    if (6'h3d == _T_253) begin
                                      mem_61 <= _GEN_20;
                                    end else begin
                                      if (6'h3d == _T_248) begin
                                        mem_61 <= _GEN_19;
                                      end else begin
                                        if (6'h3d == _T_243) begin
                                          mem_61 <= _GEN_18;
                                        end else begin
                                          if (6'h3d == _T_238) begin
                                            mem_61 <= _GEN_17;
                                          end else begin
                                            if (6'h3d == _T_233) begin
                                              mem_61 <= _GEN_16;
                                            end else begin
                                              if (6'h3d == _T_228) begin
                                                mem_61 <= _GEN_15;
                                              end else begin
                                                if (6'h3d == _T_223) begin
                                                  mem_61 <= _GEN_14;
                                                end else begin
                                                  if (6'h3d == _T_218) begin
                                                    mem_61 <= _GEN_13;
                                                  end else begin
                                                    if (6'h3d == _T_213) begin
                                                      mem_61 <= _GEN_12;
                                                    end else begin
                                                      if (6'h3d == _T_208) begin
                                                        mem_61 <= _GEN_11;
                                                      end else begin
                                                        if (6'h3d == _T_203) begin
                                                          mem_61 <= _GEN_10;
                                                        end else begin
                                                          if (6'h3d == _T_198) begin
                                                            mem_61 <= _GEN_9;
                                                          end else begin
                                                            if (6'h3d == _T_193) begin
                                                              mem_61 <= _GEN_8;
                                                            end else begin
                                                              if (6'h3d == _T_188) begin
                                                                mem_61 <= _GEN_7;
                                                              end else begin
                                                                if (6'h3d == _T_183) begin
                                                                  mem_61 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h3d == _T_178) begin
                                                                    mem_61 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h3d == _T_173) begin
                                                                      mem_61 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h3d == _T_168) begin
                                                                        mem_61 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h3d == _T_163) begin
                                                                          mem_61 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h3d == _T_158) begin
                                                                            mem_61 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h3d == _T_153) begin
                                                                              mem_61 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h3d == _T_308) begin
              mem_61 <= _GEN_31;
            end else begin
              if (6'h3d == _T_303) begin
                mem_61 <= _GEN_30;
              end else begin
                if (6'h3d == _T_298) begin
                  mem_61 <= _GEN_29;
                end else begin
                  if (6'h3d == _T_293) begin
                    mem_61 <= _GEN_28;
                  end else begin
                    if (6'h3d == _T_288) begin
                      mem_61 <= _GEN_27;
                    end else begin
                      if (6'h3d == _T_283) begin
                        mem_61 <= _GEN_26;
                      end else begin
                        if (6'h3d == _T_278) begin
                          mem_61 <= _GEN_25;
                        end else begin
                          if (6'h3d == _T_273) begin
                            mem_61 <= _GEN_24;
                          end else begin
                            if (6'h3d == _T_268) begin
                              mem_61 <= _GEN_23;
                            end else begin
                              if (6'h3d == _T_263) begin
                                mem_61 <= _GEN_22;
                              end else begin
                                if (6'h3d == _T_258) begin
                                  mem_61 <= _GEN_21;
                                end else begin
                                  if (6'h3d == _T_253) begin
                                    mem_61 <= _GEN_20;
                                  end else begin
                                    if (6'h3d == _T_248) begin
                                      mem_61 <= _GEN_19;
                                    end else begin
                                      if (6'h3d == _T_243) begin
                                        mem_61 <= _GEN_18;
                                      end else begin
                                        if (6'h3d == _T_238) begin
                                          mem_61 <= _GEN_17;
                                        end else begin
                                          if (6'h3d == _T_233) begin
                                            mem_61 <= _GEN_16;
                                          end else begin
                                            if (6'h3d == _T_228) begin
                                              mem_61 <= _GEN_15;
                                            end else begin
                                              if (6'h3d == _T_223) begin
                                                mem_61 <= _GEN_14;
                                              end else begin
                                                if (6'h3d == _T_218) begin
                                                  mem_61 <= _GEN_13;
                                                end else begin
                                                  if (6'h3d == _T_213) begin
                                                    mem_61 <= _GEN_12;
                                                  end else begin
                                                    if (6'h3d == _T_208) begin
                                                      mem_61 <= _GEN_11;
                                                    end else begin
                                                      if (6'h3d == _T_203) begin
                                                        mem_61 <= _GEN_10;
                                                      end else begin
                                                        if (6'h3d == _T_198) begin
                                                          mem_61 <= _GEN_9;
                                                        end else begin
                                                          if (6'h3d == _T_193) begin
                                                            mem_61 <= _GEN_8;
                                                          end else begin
                                                            if (6'h3d == _T_188) begin
                                                              mem_61 <= _GEN_7;
                                                            end else begin
                                                              if (6'h3d == _T_183) begin
                                                                mem_61 <= _GEN_6;
                                                              end else begin
                                                                if (6'h3d == _T_178) begin
                                                                  mem_61 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h3d == _T_173) begin
                                                                    mem_61 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h3d == _T_168) begin
                                                                      mem_61 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h3d == _T_163) begin
                                                                        mem_61 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h3d == _T_158) begin
                                                                          mem_61 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h3d == _T_153) begin
                                                                            mem_61 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h3d == _T_308) begin
            mem_61 <= _GEN_31;
          end else begin
            if (6'h3d == _T_303) begin
              mem_61 <= _GEN_30;
            end else begin
              if (6'h3d == _T_298) begin
                mem_61 <= _GEN_29;
              end else begin
                if (6'h3d == _T_293) begin
                  mem_61 <= _GEN_28;
                end else begin
                  if (6'h3d == _T_288) begin
                    mem_61 <= _GEN_27;
                  end else begin
                    if (6'h3d == _T_283) begin
                      mem_61 <= _GEN_26;
                    end else begin
                      if (6'h3d == _T_278) begin
                        mem_61 <= _GEN_25;
                      end else begin
                        if (6'h3d == _T_273) begin
                          mem_61 <= _GEN_24;
                        end else begin
                          if (6'h3d == _T_268) begin
                            mem_61 <= _GEN_23;
                          end else begin
                            if (6'h3d == _T_263) begin
                              mem_61 <= _GEN_22;
                            end else begin
                              if (6'h3d == _T_258) begin
                                mem_61 <= _GEN_21;
                              end else begin
                                if (6'h3d == _T_253) begin
                                  mem_61 <= _GEN_20;
                                end else begin
                                  if (6'h3d == _T_248) begin
                                    mem_61 <= _GEN_19;
                                  end else begin
                                    if (6'h3d == _T_243) begin
                                      mem_61 <= _GEN_18;
                                    end else begin
                                      if (6'h3d == _T_238) begin
                                        mem_61 <= _GEN_17;
                                      end else begin
                                        if (6'h3d == _T_233) begin
                                          mem_61 <= _GEN_16;
                                        end else begin
                                          if (6'h3d == _T_228) begin
                                            mem_61 <= _GEN_15;
                                          end else begin
                                            if (6'h3d == _T_223) begin
                                              mem_61 <= _GEN_14;
                                            end else begin
                                              if (6'h3d == _T_218) begin
                                                mem_61 <= _GEN_13;
                                              end else begin
                                                if (6'h3d == _T_213) begin
                                                  mem_61 <= _GEN_12;
                                                end else begin
                                                  if (6'h3d == _T_208) begin
                                                    mem_61 <= _GEN_11;
                                                  end else begin
                                                    if (6'h3d == _T_203) begin
                                                      mem_61 <= _GEN_10;
                                                    end else begin
                                                      if (6'h3d == _T_198) begin
                                                        mem_61 <= _GEN_9;
                                                      end else begin
                                                        if (6'h3d == _T_193) begin
                                                          mem_61 <= _GEN_8;
                                                        end else begin
                                                          if (6'h3d == _T_188) begin
                                                            mem_61 <= _GEN_7;
                                                          end else begin
                                                            if (6'h3d == _T_183) begin
                                                              mem_61 <= _GEN_6;
                                                            end else begin
                                                              if (6'h3d == _T_178) begin
                                                                mem_61 <= _GEN_5;
                                                              end else begin
                                                                if (6'h3d == _T_173) begin
                                                                  mem_61 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h3d == _T_168) begin
                                                                    mem_61 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h3d == _T_163) begin
                                                                      mem_61 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h3d == _T_158) begin
                                                                        mem_61 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h3d == _T_153) begin
                                                                          mem_61 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h3d == _T_308) begin
          mem_61 <= _GEN_31;
        end else begin
          if (6'h3d == _T_303) begin
            mem_61 <= _GEN_30;
          end else begin
            if (6'h3d == _T_298) begin
              mem_61 <= _GEN_29;
            end else begin
              if (6'h3d == _T_293) begin
                mem_61 <= _GEN_28;
              end else begin
                if (6'h3d == _T_288) begin
                  mem_61 <= _GEN_27;
                end else begin
                  if (6'h3d == _T_283) begin
                    mem_61 <= _GEN_26;
                  end else begin
                    if (6'h3d == _T_278) begin
                      mem_61 <= _GEN_25;
                    end else begin
                      if (6'h3d == _T_273) begin
                        mem_61 <= _GEN_24;
                      end else begin
                        if (6'h3d == _T_268) begin
                          mem_61 <= _GEN_23;
                        end else begin
                          if (6'h3d == _T_263) begin
                            mem_61 <= _GEN_22;
                          end else begin
                            if (6'h3d == _T_258) begin
                              mem_61 <= _GEN_21;
                            end else begin
                              if (6'h3d == _T_253) begin
                                mem_61 <= _GEN_20;
                              end else begin
                                if (6'h3d == _T_248) begin
                                  mem_61 <= _GEN_19;
                                end else begin
                                  if (6'h3d == _T_243) begin
                                    mem_61 <= _GEN_18;
                                  end else begin
                                    if (6'h3d == _T_238) begin
                                      mem_61 <= _GEN_17;
                                    end else begin
                                      if (6'h3d == _T_233) begin
                                        mem_61 <= _GEN_16;
                                      end else begin
                                        if (6'h3d == _T_228) begin
                                          mem_61 <= _GEN_15;
                                        end else begin
                                          if (6'h3d == _T_223) begin
                                            mem_61 <= _GEN_14;
                                          end else begin
                                            if (6'h3d == _T_218) begin
                                              mem_61 <= _GEN_13;
                                            end else begin
                                              if (6'h3d == _T_213) begin
                                                mem_61 <= _GEN_12;
                                              end else begin
                                                if (6'h3d == _T_208) begin
                                                  mem_61 <= _GEN_11;
                                                end else begin
                                                  if (6'h3d == _T_203) begin
                                                    mem_61 <= _GEN_10;
                                                  end else begin
                                                    if (6'h3d == _T_198) begin
                                                      mem_61 <= _GEN_9;
                                                    end else begin
                                                      if (6'h3d == _T_193) begin
                                                        mem_61 <= _GEN_8;
                                                      end else begin
                                                        if (6'h3d == _T_188) begin
                                                          mem_61 <= _GEN_7;
                                                        end else begin
                                                          if (6'h3d == _T_183) begin
                                                            mem_61 <= _GEN_6;
                                                          end else begin
                                                            if (6'h3d == _T_178) begin
                                                              mem_61 <= _GEN_5;
                                                            end else begin
                                                              if (6'h3d == _T_173) begin
                                                                mem_61 <= _GEN_4;
                                                              end else begin
                                                                if (6'h3d == _T_168) begin
                                                                  mem_61 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h3d == _T_163) begin
                                                                    mem_61 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h3d == _T_158) begin
                                                                      mem_61 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h3d == _T_153) begin
                                                                        mem_61 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h3e == wPos) begin
            mem_62 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h3e == _T_308) begin
                mem_62 <= _GEN_31;
              end else begin
                if (6'h3e == _T_303) begin
                  mem_62 <= _GEN_30;
                end else begin
                  if (6'h3e == _T_298) begin
                    mem_62 <= _GEN_29;
                  end else begin
                    if (6'h3e == _T_293) begin
                      mem_62 <= _GEN_28;
                    end else begin
                      if (6'h3e == _T_288) begin
                        mem_62 <= _GEN_27;
                      end else begin
                        if (6'h3e == _T_283) begin
                          mem_62 <= _GEN_26;
                        end else begin
                          if (6'h3e == _T_278) begin
                            mem_62 <= _GEN_25;
                          end else begin
                            if (6'h3e == _T_273) begin
                              mem_62 <= _GEN_24;
                            end else begin
                              if (6'h3e == _T_268) begin
                                mem_62 <= _GEN_23;
                              end else begin
                                if (6'h3e == _T_263) begin
                                  mem_62 <= _GEN_22;
                                end else begin
                                  if (6'h3e == _T_258) begin
                                    mem_62 <= _GEN_21;
                                  end else begin
                                    if (6'h3e == _T_253) begin
                                      mem_62 <= _GEN_20;
                                    end else begin
                                      if (6'h3e == _T_248) begin
                                        mem_62 <= _GEN_19;
                                      end else begin
                                        if (6'h3e == _T_243) begin
                                          mem_62 <= _GEN_18;
                                        end else begin
                                          if (6'h3e == _T_238) begin
                                            mem_62 <= _GEN_17;
                                          end else begin
                                            if (6'h3e == _T_233) begin
                                              mem_62 <= _GEN_16;
                                            end else begin
                                              if (6'h3e == _T_228) begin
                                                mem_62 <= _GEN_15;
                                              end else begin
                                                if (6'h3e == _T_223) begin
                                                  mem_62 <= _GEN_14;
                                                end else begin
                                                  if (6'h3e == _T_218) begin
                                                    mem_62 <= _GEN_13;
                                                  end else begin
                                                    if (6'h3e == _T_213) begin
                                                      mem_62 <= _GEN_12;
                                                    end else begin
                                                      if (6'h3e == _T_208) begin
                                                        mem_62 <= _GEN_11;
                                                      end else begin
                                                        if (6'h3e == _T_203) begin
                                                          mem_62 <= _GEN_10;
                                                        end else begin
                                                          if (6'h3e == _T_198) begin
                                                            mem_62 <= _GEN_9;
                                                          end else begin
                                                            if (6'h3e == _T_193) begin
                                                              mem_62 <= _GEN_8;
                                                            end else begin
                                                              if (6'h3e == _T_188) begin
                                                                mem_62 <= _GEN_7;
                                                              end else begin
                                                                if (6'h3e == _T_183) begin
                                                                  mem_62 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h3e == _T_178) begin
                                                                    mem_62 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h3e == _T_173) begin
                                                                      mem_62 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h3e == _T_168) begin
                                                                        mem_62 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h3e == _T_163) begin
                                                                          mem_62 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h3e == _T_158) begin
                                                                            mem_62 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h3e == _T_153) begin
                                                                              mem_62 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h3e == _T_308) begin
              mem_62 <= _GEN_31;
            end else begin
              if (6'h3e == _T_303) begin
                mem_62 <= _GEN_30;
              end else begin
                if (6'h3e == _T_298) begin
                  mem_62 <= _GEN_29;
                end else begin
                  if (6'h3e == _T_293) begin
                    mem_62 <= _GEN_28;
                  end else begin
                    if (6'h3e == _T_288) begin
                      mem_62 <= _GEN_27;
                    end else begin
                      if (6'h3e == _T_283) begin
                        mem_62 <= _GEN_26;
                      end else begin
                        if (6'h3e == _T_278) begin
                          mem_62 <= _GEN_25;
                        end else begin
                          if (6'h3e == _T_273) begin
                            mem_62 <= _GEN_24;
                          end else begin
                            if (6'h3e == _T_268) begin
                              mem_62 <= _GEN_23;
                            end else begin
                              if (6'h3e == _T_263) begin
                                mem_62 <= _GEN_22;
                              end else begin
                                if (6'h3e == _T_258) begin
                                  mem_62 <= _GEN_21;
                                end else begin
                                  if (6'h3e == _T_253) begin
                                    mem_62 <= _GEN_20;
                                  end else begin
                                    if (6'h3e == _T_248) begin
                                      mem_62 <= _GEN_19;
                                    end else begin
                                      if (6'h3e == _T_243) begin
                                        mem_62 <= _GEN_18;
                                      end else begin
                                        if (6'h3e == _T_238) begin
                                          mem_62 <= _GEN_17;
                                        end else begin
                                          if (6'h3e == _T_233) begin
                                            mem_62 <= _GEN_16;
                                          end else begin
                                            if (6'h3e == _T_228) begin
                                              mem_62 <= _GEN_15;
                                            end else begin
                                              if (6'h3e == _T_223) begin
                                                mem_62 <= _GEN_14;
                                              end else begin
                                                if (6'h3e == _T_218) begin
                                                  mem_62 <= _GEN_13;
                                                end else begin
                                                  if (6'h3e == _T_213) begin
                                                    mem_62 <= _GEN_12;
                                                  end else begin
                                                    if (6'h3e == _T_208) begin
                                                      mem_62 <= _GEN_11;
                                                    end else begin
                                                      if (6'h3e == _T_203) begin
                                                        mem_62 <= _GEN_10;
                                                      end else begin
                                                        if (6'h3e == _T_198) begin
                                                          mem_62 <= _GEN_9;
                                                        end else begin
                                                          if (6'h3e == _T_193) begin
                                                            mem_62 <= _GEN_8;
                                                          end else begin
                                                            if (6'h3e == _T_188) begin
                                                              mem_62 <= _GEN_7;
                                                            end else begin
                                                              if (6'h3e == _T_183) begin
                                                                mem_62 <= _GEN_6;
                                                              end else begin
                                                                if (6'h3e == _T_178) begin
                                                                  mem_62 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h3e == _T_173) begin
                                                                    mem_62 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h3e == _T_168) begin
                                                                      mem_62 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h3e == _T_163) begin
                                                                        mem_62 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h3e == _T_158) begin
                                                                          mem_62 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h3e == _T_153) begin
                                                                            mem_62 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h3e == _T_308) begin
            mem_62 <= _GEN_31;
          end else begin
            if (6'h3e == _T_303) begin
              mem_62 <= _GEN_30;
            end else begin
              if (6'h3e == _T_298) begin
                mem_62 <= _GEN_29;
              end else begin
                if (6'h3e == _T_293) begin
                  mem_62 <= _GEN_28;
                end else begin
                  if (6'h3e == _T_288) begin
                    mem_62 <= _GEN_27;
                  end else begin
                    if (6'h3e == _T_283) begin
                      mem_62 <= _GEN_26;
                    end else begin
                      if (6'h3e == _T_278) begin
                        mem_62 <= _GEN_25;
                      end else begin
                        if (6'h3e == _T_273) begin
                          mem_62 <= _GEN_24;
                        end else begin
                          if (6'h3e == _T_268) begin
                            mem_62 <= _GEN_23;
                          end else begin
                            if (6'h3e == _T_263) begin
                              mem_62 <= _GEN_22;
                            end else begin
                              if (6'h3e == _T_258) begin
                                mem_62 <= _GEN_21;
                              end else begin
                                if (6'h3e == _T_253) begin
                                  mem_62 <= _GEN_20;
                                end else begin
                                  if (6'h3e == _T_248) begin
                                    mem_62 <= _GEN_19;
                                  end else begin
                                    if (6'h3e == _T_243) begin
                                      mem_62 <= _GEN_18;
                                    end else begin
                                      if (6'h3e == _T_238) begin
                                        mem_62 <= _GEN_17;
                                      end else begin
                                        if (6'h3e == _T_233) begin
                                          mem_62 <= _GEN_16;
                                        end else begin
                                          if (6'h3e == _T_228) begin
                                            mem_62 <= _GEN_15;
                                          end else begin
                                            if (6'h3e == _T_223) begin
                                              mem_62 <= _GEN_14;
                                            end else begin
                                              if (6'h3e == _T_218) begin
                                                mem_62 <= _GEN_13;
                                              end else begin
                                                if (6'h3e == _T_213) begin
                                                  mem_62 <= _GEN_12;
                                                end else begin
                                                  if (6'h3e == _T_208) begin
                                                    mem_62 <= _GEN_11;
                                                  end else begin
                                                    if (6'h3e == _T_203) begin
                                                      mem_62 <= _GEN_10;
                                                    end else begin
                                                      if (6'h3e == _T_198) begin
                                                        mem_62 <= _GEN_9;
                                                      end else begin
                                                        if (6'h3e == _T_193) begin
                                                          mem_62 <= _GEN_8;
                                                        end else begin
                                                          if (6'h3e == _T_188) begin
                                                            mem_62 <= _GEN_7;
                                                          end else begin
                                                            if (6'h3e == _T_183) begin
                                                              mem_62 <= _GEN_6;
                                                            end else begin
                                                              if (6'h3e == _T_178) begin
                                                                mem_62 <= _GEN_5;
                                                              end else begin
                                                                if (6'h3e == _T_173) begin
                                                                  mem_62 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h3e == _T_168) begin
                                                                    mem_62 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h3e == _T_163) begin
                                                                      mem_62 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h3e == _T_158) begin
                                                                        mem_62 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h3e == _T_153) begin
                                                                          mem_62 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h3e == _T_308) begin
          mem_62 <= _GEN_31;
        end else begin
          if (6'h3e == _T_303) begin
            mem_62 <= _GEN_30;
          end else begin
            if (6'h3e == _T_298) begin
              mem_62 <= _GEN_29;
            end else begin
              if (6'h3e == _T_293) begin
                mem_62 <= _GEN_28;
              end else begin
                if (6'h3e == _T_288) begin
                  mem_62 <= _GEN_27;
                end else begin
                  if (6'h3e == _T_283) begin
                    mem_62 <= _GEN_26;
                  end else begin
                    if (6'h3e == _T_278) begin
                      mem_62 <= _GEN_25;
                    end else begin
                      if (6'h3e == _T_273) begin
                        mem_62 <= _GEN_24;
                      end else begin
                        if (6'h3e == _T_268) begin
                          mem_62 <= _GEN_23;
                        end else begin
                          if (6'h3e == _T_263) begin
                            mem_62 <= _GEN_22;
                          end else begin
                            if (6'h3e == _T_258) begin
                              mem_62 <= _GEN_21;
                            end else begin
                              if (6'h3e == _T_253) begin
                                mem_62 <= _GEN_20;
                              end else begin
                                if (6'h3e == _T_248) begin
                                  mem_62 <= _GEN_19;
                                end else begin
                                  if (6'h3e == _T_243) begin
                                    mem_62 <= _GEN_18;
                                  end else begin
                                    if (6'h3e == _T_238) begin
                                      mem_62 <= _GEN_17;
                                    end else begin
                                      if (6'h3e == _T_233) begin
                                        mem_62 <= _GEN_16;
                                      end else begin
                                        if (6'h3e == _T_228) begin
                                          mem_62 <= _GEN_15;
                                        end else begin
                                          if (6'h3e == _T_223) begin
                                            mem_62 <= _GEN_14;
                                          end else begin
                                            if (6'h3e == _T_218) begin
                                              mem_62 <= _GEN_13;
                                            end else begin
                                              if (6'h3e == _T_213) begin
                                                mem_62 <= _GEN_12;
                                              end else begin
                                                if (6'h3e == _T_208) begin
                                                  mem_62 <= _GEN_11;
                                                end else begin
                                                  if (6'h3e == _T_203) begin
                                                    mem_62 <= _GEN_10;
                                                  end else begin
                                                    if (6'h3e == _T_198) begin
                                                      mem_62 <= _GEN_9;
                                                    end else begin
                                                      if (6'h3e == _T_193) begin
                                                        mem_62 <= _GEN_8;
                                                      end else begin
                                                        if (6'h3e == _T_188) begin
                                                          mem_62 <= _GEN_7;
                                                        end else begin
                                                          if (6'h3e == _T_183) begin
                                                            mem_62 <= _GEN_6;
                                                          end else begin
                                                            if (6'h3e == _T_178) begin
                                                              mem_62 <= _GEN_5;
                                                            end else begin
                                                              if (6'h3e == _T_173) begin
                                                                mem_62 <= _GEN_4;
                                                              end else begin
                                                                if (6'h3e == _T_168) begin
                                                                  mem_62 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h3e == _T_163) begin
                                                                    mem_62 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h3e == _T_158) begin
                                                                      mem_62 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h3e == _T_153) begin
                                                                        mem_62 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_315) begin
      if (io_push) begin
        if (_T_149) begin
          if (6'h3f == wPos) begin
            mem_63 <= _GEN_32;
          end else begin
            if (_T_150) begin
              if (6'h3f == _T_308) begin
                mem_63 <= _GEN_31;
              end else begin
                if (6'h3f == _T_303) begin
                  mem_63 <= _GEN_30;
                end else begin
                  if (6'h3f == _T_298) begin
                    mem_63 <= _GEN_29;
                  end else begin
                    if (6'h3f == _T_293) begin
                      mem_63 <= _GEN_28;
                    end else begin
                      if (6'h3f == _T_288) begin
                        mem_63 <= _GEN_27;
                      end else begin
                        if (6'h3f == _T_283) begin
                          mem_63 <= _GEN_26;
                        end else begin
                          if (6'h3f == _T_278) begin
                            mem_63 <= _GEN_25;
                          end else begin
                            if (6'h3f == _T_273) begin
                              mem_63 <= _GEN_24;
                            end else begin
                              if (6'h3f == _T_268) begin
                                mem_63 <= _GEN_23;
                              end else begin
                                if (6'h3f == _T_263) begin
                                  mem_63 <= _GEN_22;
                                end else begin
                                  if (6'h3f == _T_258) begin
                                    mem_63 <= _GEN_21;
                                  end else begin
                                    if (6'h3f == _T_253) begin
                                      mem_63 <= _GEN_20;
                                    end else begin
                                      if (6'h3f == _T_248) begin
                                        mem_63 <= _GEN_19;
                                      end else begin
                                        if (6'h3f == _T_243) begin
                                          mem_63 <= _GEN_18;
                                        end else begin
                                          if (6'h3f == _T_238) begin
                                            mem_63 <= _GEN_17;
                                          end else begin
                                            if (6'h3f == _T_233) begin
                                              mem_63 <= _GEN_16;
                                            end else begin
                                              if (6'h3f == _T_228) begin
                                                mem_63 <= _GEN_15;
                                              end else begin
                                                if (6'h3f == _T_223) begin
                                                  mem_63 <= _GEN_14;
                                                end else begin
                                                  if (6'h3f == _T_218) begin
                                                    mem_63 <= _GEN_13;
                                                  end else begin
                                                    if (6'h3f == _T_213) begin
                                                      mem_63 <= _GEN_12;
                                                    end else begin
                                                      if (6'h3f == _T_208) begin
                                                        mem_63 <= _GEN_11;
                                                      end else begin
                                                        if (6'h3f == _T_203) begin
                                                          mem_63 <= _GEN_10;
                                                        end else begin
                                                          if (6'h3f == _T_198) begin
                                                            mem_63 <= _GEN_9;
                                                          end else begin
                                                            if (6'h3f == _T_193) begin
                                                              mem_63 <= _GEN_8;
                                                            end else begin
                                                              if (6'h3f == _T_188) begin
                                                                mem_63 <= _GEN_7;
                                                              end else begin
                                                                if (6'h3f == _T_183) begin
                                                                  mem_63 <= _GEN_6;
                                                                end else begin
                                                                  if (6'h3f == _T_178) begin
                                                                    mem_63 <= _GEN_5;
                                                                  end else begin
                                                                    if (6'h3f == _T_173) begin
                                                                      mem_63 <= _GEN_4;
                                                                    end else begin
                                                                      if (6'h3f == _T_168) begin
                                                                        mem_63 <= _GEN_3;
                                                                      end else begin
                                                                        if (6'h3f == _T_163) begin
                                                                          mem_63 <= _GEN_2;
                                                                        end else begin
                                                                          if (6'h3f == _T_158) begin
                                                                            mem_63 <= _GEN_1;
                                                                          end else begin
                                                                            if (6'h3f == _T_153) begin
                                                                              mem_63 <= _GEN_0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_150) begin
            if (6'h3f == _T_308) begin
              mem_63 <= _GEN_31;
            end else begin
              if (6'h3f == _T_303) begin
                mem_63 <= _GEN_30;
              end else begin
                if (6'h3f == _T_298) begin
                  mem_63 <= _GEN_29;
                end else begin
                  if (6'h3f == _T_293) begin
                    mem_63 <= _GEN_28;
                  end else begin
                    if (6'h3f == _T_288) begin
                      mem_63 <= _GEN_27;
                    end else begin
                      if (6'h3f == _T_283) begin
                        mem_63 <= _GEN_26;
                      end else begin
                        if (6'h3f == _T_278) begin
                          mem_63 <= _GEN_25;
                        end else begin
                          if (6'h3f == _T_273) begin
                            mem_63 <= _GEN_24;
                          end else begin
                            if (6'h3f == _T_268) begin
                              mem_63 <= _GEN_23;
                            end else begin
                              if (6'h3f == _T_263) begin
                                mem_63 <= _GEN_22;
                              end else begin
                                if (6'h3f == _T_258) begin
                                  mem_63 <= _GEN_21;
                                end else begin
                                  if (6'h3f == _T_253) begin
                                    mem_63 <= _GEN_20;
                                  end else begin
                                    if (6'h3f == _T_248) begin
                                      mem_63 <= _GEN_19;
                                    end else begin
                                      if (6'h3f == _T_243) begin
                                        mem_63 <= _GEN_18;
                                      end else begin
                                        if (6'h3f == _T_238) begin
                                          mem_63 <= _GEN_17;
                                        end else begin
                                          if (6'h3f == _T_233) begin
                                            mem_63 <= _GEN_16;
                                          end else begin
                                            if (6'h3f == _T_228) begin
                                              mem_63 <= _GEN_15;
                                            end else begin
                                              if (6'h3f == _T_223) begin
                                                mem_63 <= _GEN_14;
                                              end else begin
                                                if (6'h3f == _T_218) begin
                                                  mem_63 <= _GEN_13;
                                                end else begin
                                                  if (6'h3f == _T_213) begin
                                                    mem_63 <= _GEN_12;
                                                  end else begin
                                                    if (6'h3f == _T_208) begin
                                                      mem_63 <= _GEN_11;
                                                    end else begin
                                                      if (6'h3f == _T_203) begin
                                                        mem_63 <= _GEN_10;
                                                      end else begin
                                                        if (6'h3f == _T_198) begin
                                                          mem_63 <= _GEN_9;
                                                        end else begin
                                                          if (6'h3f == _T_193) begin
                                                            mem_63 <= _GEN_8;
                                                          end else begin
                                                            if (6'h3f == _T_188) begin
                                                              mem_63 <= _GEN_7;
                                                            end else begin
                                                              if (6'h3f == _T_183) begin
                                                                mem_63 <= _GEN_6;
                                                              end else begin
                                                                if (6'h3f == _T_178) begin
                                                                  mem_63 <= _GEN_5;
                                                                end else begin
                                                                  if (6'h3f == _T_173) begin
                                                                    mem_63 <= _GEN_4;
                                                                  end else begin
                                                                    if (6'h3f == _T_168) begin
                                                                      mem_63 <= _GEN_3;
                                                                    end else begin
                                                                      if (6'h3f == _T_163) begin
                                                                        mem_63 <= _GEN_2;
                                                                      end else begin
                                                                        if (6'h3f == _T_158) begin
                                                                          mem_63 <= _GEN_1;
                                                                        end else begin
                                                                          if (6'h3f == _T_153) begin
                                                                            mem_63 <= _GEN_0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_150) begin
          if (6'h3f == _T_308) begin
            mem_63 <= _GEN_31;
          end else begin
            if (6'h3f == _T_303) begin
              mem_63 <= _GEN_30;
            end else begin
              if (6'h3f == _T_298) begin
                mem_63 <= _GEN_29;
              end else begin
                if (6'h3f == _T_293) begin
                  mem_63 <= _GEN_28;
                end else begin
                  if (6'h3f == _T_288) begin
                    mem_63 <= _GEN_27;
                  end else begin
                    if (6'h3f == _T_283) begin
                      mem_63 <= _GEN_26;
                    end else begin
                      if (6'h3f == _T_278) begin
                        mem_63 <= _GEN_25;
                      end else begin
                        if (6'h3f == _T_273) begin
                          mem_63 <= _GEN_24;
                        end else begin
                          if (6'h3f == _T_268) begin
                            mem_63 <= _GEN_23;
                          end else begin
                            if (6'h3f == _T_263) begin
                              mem_63 <= _GEN_22;
                            end else begin
                              if (6'h3f == _T_258) begin
                                mem_63 <= _GEN_21;
                              end else begin
                                if (6'h3f == _T_253) begin
                                  mem_63 <= _GEN_20;
                                end else begin
                                  if (6'h3f == _T_248) begin
                                    mem_63 <= _GEN_19;
                                  end else begin
                                    if (6'h3f == _T_243) begin
                                      mem_63 <= _GEN_18;
                                    end else begin
                                      if (6'h3f == _T_238) begin
                                        mem_63 <= _GEN_17;
                                      end else begin
                                        if (6'h3f == _T_233) begin
                                          mem_63 <= _GEN_16;
                                        end else begin
                                          if (6'h3f == _T_228) begin
                                            mem_63 <= _GEN_15;
                                          end else begin
                                            if (6'h3f == _T_223) begin
                                              mem_63 <= _GEN_14;
                                            end else begin
                                              if (6'h3f == _T_218) begin
                                                mem_63 <= _GEN_13;
                                              end else begin
                                                if (6'h3f == _T_213) begin
                                                  mem_63 <= _GEN_12;
                                                end else begin
                                                  if (6'h3f == _T_208) begin
                                                    mem_63 <= _GEN_11;
                                                  end else begin
                                                    if (6'h3f == _T_203) begin
                                                      mem_63 <= _GEN_10;
                                                    end else begin
                                                      if (6'h3f == _T_198) begin
                                                        mem_63 <= _GEN_9;
                                                      end else begin
                                                        if (6'h3f == _T_193) begin
                                                          mem_63 <= _GEN_8;
                                                        end else begin
                                                          if (6'h3f == _T_188) begin
                                                            mem_63 <= _GEN_7;
                                                          end else begin
                                                            if (6'h3f == _T_183) begin
                                                              mem_63 <= _GEN_6;
                                                            end else begin
                                                              if (6'h3f == _T_178) begin
                                                                mem_63 <= _GEN_5;
                                                              end else begin
                                                                if (6'h3f == _T_173) begin
                                                                  mem_63 <= _GEN_4;
                                                                end else begin
                                                                  if (6'h3f == _T_168) begin
                                                                    mem_63 <= _GEN_3;
                                                                  end else begin
                                                                    if (6'h3f == _T_163) begin
                                                                      mem_63 <= _GEN_2;
                                                                    end else begin
                                                                      if (6'h3f == _T_158) begin
                                                                        mem_63 <= _GEN_1;
                                                                      end else begin
                                                                        if (6'h3f == _T_153) begin
                                                                          mem_63 <= _GEN_0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_150) begin
        if (6'h3f == _T_308) begin
          mem_63 <= _GEN_31;
        end else begin
          if (6'h3f == _T_303) begin
            mem_63 <= _GEN_30;
          end else begin
            if (6'h3f == _T_298) begin
              mem_63 <= _GEN_29;
            end else begin
              if (6'h3f == _T_293) begin
                mem_63 <= _GEN_28;
              end else begin
                if (6'h3f == _T_288) begin
                  mem_63 <= _GEN_27;
                end else begin
                  if (6'h3f == _T_283) begin
                    mem_63 <= _GEN_26;
                  end else begin
                    if (6'h3f == _T_278) begin
                      mem_63 <= _GEN_25;
                    end else begin
                      if (6'h3f == _T_273) begin
                        mem_63 <= _GEN_24;
                      end else begin
                        if (6'h3f == _T_268) begin
                          mem_63 <= _GEN_23;
                        end else begin
                          if (6'h3f == _T_263) begin
                            mem_63 <= _GEN_22;
                          end else begin
                            if (6'h3f == _T_258) begin
                              mem_63 <= _GEN_21;
                            end else begin
                              if (6'h3f == _T_253) begin
                                mem_63 <= _GEN_20;
                              end else begin
                                if (6'h3f == _T_248) begin
                                  mem_63 <= _GEN_19;
                                end else begin
                                  if (6'h3f == _T_243) begin
                                    mem_63 <= _GEN_18;
                                  end else begin
                                    if (6'h3f == _T_238) begin
                                      mem_63 <= _GEN_17;
                                    end else begin
                                      if (6'h3f == _T_233) begin
                                        mem_63 <= _GEN_16;
                                      end else begin
                                        if (6'h3f == _T_228) begin
                                          mem_63 <= _GEN_15;
                                        end else begin
                                          if (6'h3f == _T_223) begin
                                            mem_63 <= _GEN_14;
                                          end else begin
                                            if (6'h3f == _T_218) begin
                                              mem_63 <= _GEN_13;
                                            end else begin
                                              if (6'h3f == _T_213) begin
                                                mem_63 <= _GEN_12;
                                              end else begin
                                                if (6'h3f == _T_208) begin
                                                  mem_63 <= _GEN_11;
                                                end else begin
                                                  if (6'h3f == _T_203) begin
                                                    mem_63 <= _GEN_10;
                                                  end else begin
                                                    if (6'h3f == _T_198) begin
                                                      mem_63 <= _GEN_9;
                                                    end else begin
                                                      if (6'h3f == _T_193) begin
                                                        mem_63 <= _GEN_8;
                                                      end else begin
                                                        if (6'h3f == _T_188) begin
                                                          mem_63 <= _GEN_7;
                                                        end else begin
                                                          if (6'h3f == _T_183) begin
                                                            mem_63 <= _GEN_6;
                                                          end else begin
                                                            if (6'h3f == _T_178) begin
                                                              mem_63 <= _GEN_5;
                                                            end else begin
                                                              if (6'h3f == _T_173) begin
                                                                mem_63 <= _GEN_4;
                                                              end else begin
                                                                if (6'h3f == _T_168) begin
                                                                  mem_63 <= _GEN_3;
                                                                end else begin
                                                                  if (6'h3f == _T_163) begin
                                                                    mem_63 <= _GEN_2;
                                                                  end else begin
                                                                    if (6'h3f == _T_158) begin
                                                                      mem_63 <= _GEN_1;
                                                                    end else begin
                                                                      if (6'h3f == _T_153) begin
                                                                        mem_63 <= _GEN_0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module XNOR(
  input  [31:0] io_in1,
  input  [31:0] io_in2_0,
  input  [31:0] io_in2_1,
  input  [31:0] io_in2_2,
  input  [31:0] io_in2_3,
  output [31:0] io_out_0,
  output [31:0] io_out_1,
  output [31:0] io_out_2,
  output [31:0] io_out_3
);
  wire [31:0] _T_21;
  wire [31:0] _T_22;
  wire [31:0] _T_23;
  wire [31:0] _T_24;
  wire [31:0] _T_25;
  wire [31:0] _T_26;
  wire [31:0] _T_27;
  wire [31:0] _T_28;
  assign io_out_0 = _T_22;
  assign io_out_1 = _T_24;
  assign io_out_2 = _T_26;
  assign io_out_3 = _T_28;
  assign _T_21 = io_in1 ^ io_in2_0;
  assign _T_22 = ~ _T_21;
  assign _T_23 = io_in1 ^ io_in2_1;
  assign _T_24 = ~ _T_23;
  assign _T_25 = io_in1 ^ io_in2_2;
  assign _T_26 = ~ _T_25;
  assign _T_27 = io_in1 ^ io_in2_3;
  assign _T_28 = ~ _T_27;
endmodule
module MeanBuffer(
  input         clock,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [15:0] io_cntInverse65536,
  input         io_reset,
  output [31:0] io_out
);
  reg [31:0] acc;
  reg [31:0] _GEN_5;
  reg [31:0] result;
  reg [31:0] _GEN_6;
  wire  _T_17;
  wire [32:0] _T_19;
  wire [31:0] _T_20;
  wire [31:0] _T_21;
  wire [31:0] _T_22;
  wire [31:0] _T_23;
  wire  _T_25;
  wire [32:0] _T_27;
  wire [31:0] _T_28;
  wire [31:0] _T_29;
  wire [31:0] _T_30;
  wire [31:0] _T_31;
  wire  _T_33;
  wire [32:0] _T_35;
  wire [31:0] _T_36;
  wire [31:0] _T_37;
  wire [31:0] _T_38;
  wire [31:0] _T_39;
  wire  _T_41;
  wire [32:0] _T_43;
  wire [31:0] _T_44;
  wire [31:0] _T_45;
  wire [31:0] _T_46;
  wire [31:0] _T_47;
  wire [32:0] _T_48;
  wire [31:0] _T_49;
  wire [32:0] _T_50;
  wire [31:0] _T_51;
  wire [32:0] _T_52;
  wire [31:0] absSum;
  wire  _T_54;
  wire [32:0] _T_55;
  wire [31:0] _T_56;
  wire [31:0] _GEN_4;
  wire [47:0] _T_59;
  wire [31:0] _T_60;
  wire [31:0] _GEN_0;
  wire [31:0] _GEN_1;
  wire  _T_62;
  wire [47:0] _T_63;
  wire [31:0] _T_64;
  wire [31:0] _GEN_2;
  wire [31:0] _GEN_3;
  assign io_out = result;
  assign _T_17 = $signed(io_in_0) > $signed(32'sh0);
  assign _T_19 = $signed(32'sh0) - $signed(io_in_0);
  assign _T_20 = _T_19[31:0];
  assign _T_21 = $signed(_T_20);
  assign _T_22 = _T_17 ? $signed(io_in_0) : $signed(_T_21);
  assign _T_23 = $unsigned(_T_22);
  assign _T_25 = $signed(io_in_1) > $signed(32'sh0);
  assign _T_27 = $signed(32'sh0) - $signed(io_in_1);
  assign _T_28 = _T_27[31:0];
  assign _T_29 = $signed(_T_28);
  assign _T_30 = _T_25 ? $signed(io_in_1) : $signed(_T_29);
  assign _T_31 = $unsigned(_T_30);
  assign _T_33 = $signed(io_in_2) > $signed(32'sh0);
  assign _T_35 = $signed(32'sh0) - $signed(io_in_2);
  assign _T_36 = _T_35[31:0];
  assign _T_37 = $signed(_T_36);
  assign _T_38 = _T_33 ? $signed(io_in_2) : $signed(_T_37);
  assign _T_39 = $unsigned(_T_38);
  assign _T_41 = $signed(io_in_3) > $signed(32'sh0);
  assign _T_43 = $signed(32'sh0) - $signed(io_in_3);
  assign _T_44 = _T_43[31:0];
  assign _T_45 = $signed(_T_44);
  assign _T_46 = _T_41 ? $signed(io_in_3) : $signed(_T_45);
  assign _T_47 = $unsigned(_T_46);
  assign _T_48 = _T_23 + _T_31;
  assign _T_49 = _T_48[31:0];
  assign _T_50 = _T_39 + _T_47;
  assign _T_51 = _T_50[31:0];
  assign _T_52 = _T_49 + _T_51;
  assign absSum = _T_52[31:0];
  assign _T_54 = io_reset == 1'h0;
  assign _T_55 = acc + absSum;
  assign _T_56 = _T_55[31:0];
  assign _GEN_4 = {{16'd0}, io_cntInverse65536};
  assign _T_59 = _T_56 * _GEN_4;
  assign _T_60 = _T_59[47:16];
  assign _GEN_0 = _T_54 ? _T_56 : acc;
  assign _GEN_1 = _T_54 ? _T_60 : result;
  assign _T_62 = _T_54 == 1'h0;
  assign _T_63 = absSum * _GEN_4;
  assign _T_64 = _T_63[47:16];
  assign _GEN_2 = _T_62 ? absSum : _GEN_0;
  assign _GEN_3 = _T_62 ? _T_64 : _GEN_1;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_5 = {1{$random}};
  acc = _GEN_5[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_6 = {1{$random}};
  result = _GEN_6[31:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (_T_62) begin
      acc <= absSum;
    end else begin
      if (_T_54) begin
        acc <= _T_56;
      end
    end
    if (_T_62) begin
      result <= _T_64;
    end else begin
      if (_T_54) begin
        result <= _T_60;
      end
    end
  end
endmodule
module DelayedOutput(
  input         clock,
  input         reset,
  input         io_reset,
  input  [31:0] io_input,
  input         io_update,
  output [31:0] io_output
);
  reg [31:0] reg$;
  reg [31:0] _GEN_2;
  wire  _T_9;
  wire [31:0] _GEN_0;
  wire  _T_11;
  wire  _T_12;
  wire [31:0] _GEN_1;
  assign io_output = reg$;
  assign _T_9 = reset == 1'h0;
  assign _GEN_0 = io_reset ? 32'h1 : reg$;
  assign _T_11 = io_reset == 1'h0;
  assign _T_12 = _T_11 & io_update;
  assign _GEN_1 = _T_12 ? io_input : _GEN_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2 = {1{$random}};
  reg$ = _GEN_2[31:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (_T_12) begin
      reg$ <= io_input;
    end else begin
      if (io_reset) begin
        reg$ <= 32'h1;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_reset & _T_9) begin
          $fwrite(32'h80000002,"Delay reset! %d\n",reg$);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_12 & _T_9) begin
          $fwrite(32'h80000002,"Delay Update! %d\n",io_input);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module MaxBuffer(
  input         clock,
  input         io_reset,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [3:0]  io_offset,
  output [3:0]  io_out,
  input  [3:0]  io_maxLen
);
  reg [3:0] idxReg;
  reg [31:0] _GEN_6;
  reg [31:0] dataReg;
  reg [31:0] _GEN_7;
  wire [4:0] _T_19;
  wire [3:0] _T_20;
  wire [4:0] _T_22;
  wire [3:0] _T_23;
  wire [4:0] _T_25;
  wire [3:0] _T_26;
  wire [4:0] _T_28;
  wire [3:0] _T_29;
  wire  _T_30;
  wire  _T_31;
  wire  _T_32;
  wire [3:0] _T_33;
  wire [31:0] _T_34;
  wire  _T_35;
  wire  _T_36;
  wire  _T_37;
  wire [3:0] _T_38;
  wire [31:0] _T_39;
  wire  _T_40;
  wire  _T_41;
  wire  _T_42;
  wire [3:0] _T_43;
  wire [31:0] _T_44;
  wire  cmp2;
  wire  _T_46;
  wire [31:0] _T_47;
  wire [3:0] _T_48;
  wire [31:0] _GEN_0;
  wire [3:0] _GEN_1;
  wire  _T_50;
  wire [31:0] _GEN_2;
  wire [3:0] _GEN_3;
  wire [31:0] _GEN_4;
  wire [3:0] _GEN_5;
  assign io_out = idxReg;
  assign _T_19 = 4'h0 + io_offset;
  assign _T_20 = _T_19[3:0];
  assign _T_22 = 4'h1 + io_offset;
  assign _T_23 = _T_22[3:0];
  assign _T_25 = 4'h2 + io_offset;
  assign _T_26 = _T_25[3:0];
  assign _T_28 = 4'h3 + io_offset;
  assign _T_29 = _T_28[3:0];
  assign _T_30 = $signed(io_in_0) > $signed(io_in_1);
  assign _T_31 = _T_23 >= io_maxLen;
  assign _T_32 = _T_30 | _T_31;
  assign _T_33 = _T_32 ? _T_20 : _T_23;
  assign _T_34 = _T_32 ? $signed(io_in_0) : $signed(io_in_1);
  assign _T_35 = $signed(io_in_2) > $signed(io_in_3);
  assign _T_36 = _T_29 >= io_maxLen;
  assign _T_37 = _T_35 | _T_36;
  assign _T_38 = _T_37 ? _T_26 : _T_29;
  assign _T_39 = _T_37 ? $signed(io_in_2) : $signed(io_in_3);
  assign _T_40 = $signed(_T_34) > $signed(_T_39);
  assign _T_41 = _T_38 >= io_maxLen;
  assign _T_42 = _T_40 | _T_41;
  assign _T_43 = _T_42 ? _T_33 : _T_38;
  assign _T_44 = _T_42 ? $signed(_T_34) : $signed(_T_39);
  assign cmp2 = $signed(dataReg) > $signed(_T_44);
  assign _T_46 = io_reset == 1'h0;
  assign _T_47 = cmp2 ? $signed(dataReg) : $signed(_T_44);
  assign _T_48 = cmp2 ? idxReg : _T_43;
  assign _GEN_0 = _T_46 ? $signed(_T_47) : $signed(dataReg);
  assign _GEN_1 = _T_46 ? _T_48 : idxReg;
  assign _T_50 = _T_46 == 1'h0;
  assign _GEN_2 = _T_50 ? $signed(_T_44) : $signed(_GEN_0);
  assign _GEN_3 = _T_50 ? _T_43 : _GEN_1;
  assign _GEN_4 = io_en ? $signed(_GEN_2) : $signed(dataReg);
  assign _GEN_5 = io_en ? _GEN_3 : idxReg;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_6 = {1{$random}};
  idxReg = _GEN_6[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_7 = {1{$random}};
  dataReg = _GEN_7[31:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (io_en) begin
      if (_T_50) begin
        if (_T_42) begin
          if (_T_32) begin
            idxReg <= _T_20;
          end else begin
            idxReg <= _T_23;
          end
        end else begin
          if (_T_37) begin
            idxReg <= _T_26;
          end else begin
            idxReg <= _T_29;
          end
        end
      end else begin
        if (_T_46) begin
          if (!(cmp2)) begin
            if (_T_42) begin
              if (_T_32) begin
                idxReg <= _T_20;
              end else begin
                idxReg <= _T_23;
              end
            end else begin
              if (_T_37) begin
                idxReg <= _T_26;
              end else begin
                idxReg <= _T_29;
              end
            end
          end
        end
      end
    end
    if (io_en) begin
      if (_T_50) begin
        if (_T_42) begin
          if (_T_32) begin
            dataReg <= io_in_0;
          end else begin
            dataReg <= io_in_1;
          end
        end else begin
          if (_T_37) begin
            dataReg <= io_in_2;
          end else begin
            dataReg <= io_in_3;
          end
        end
      end else begin
        if (_T_46) begin
          if (!(cmp2)) begin
            if (_T_42) begin
              if (_T_32) begin
                dataReg <= io_in_0;
              end else begin
                dataReg <= io_in_1;
              end
            end else begin
              if (_T_37) begin
                dataReg <= io_in_2;
              end else begin
                dataReg <= io_in_3;
              end
            end
          end
        end
      end
    end
  end
endmodule
module Accumulator(
  input        clock,
  input        reset,
  input  [9:0] io_in,
  output [9:0] io_out,
  input  [4:0] io_sel,
  input        io_en,
  input        io_reset
);
  reg [9:0] accumulator_0;
  reg [31:0] _GEN_131;
  reg [9:0] accumulator_1;
  reg [31:0] _GEN_132;
  reg [9:0] accumulator_2;
  reg [31:0] _GEN_133;
  reg [9:0] accumulator_3;
  reg [31:0] _GEN_134;
  reg [9:0] accumulator_4;
  reg [31:0] _GEN_135;
  reg [9:0] accumulator_5;
  reg [31:0] _GEN_136;
  reg [9:0] accumulator_6;
  reg [31:0] _GEN_137;
  reg [9:0] accumulator_7;
  reg [31:0] _GEN_138;
  reg [9:0] accumulator_8;
  reg [31:0] _GEN_139;
  reg [9:0] accumulator_9;
  reg [31:0] _GEN_140;
  reg [9:0] accumulator_10;
  reg [31:0] _GEN_141;
  reg [9:0] accumulator_11;
  reg [31:0] _GEN_142;
  reg [9:0] accumulator_12;
  reg [31:0] _GEN_143;
  reg [9:0] accumulator_13;
  reg [31:0] _GEN_144;
  reg [9:0] accumulator_14;
  reg [31:0] _GEN_145;
  reg [9:0] accumulator_15;
  reg [31:0] _GEN_146;
  reg [9:0] accumulator_16;
  reg [31:0] _GEN_147;
  reg [9:0] accumulator_17;
  reg [31:0] _GEN_148;
  reg [9:0] accumulator_18;
  reg [31:0] _GEN_149;
  reg [9:0] accumulator_19;
  reg [31:0] _GEN_150;
  reg [9:0] accumulator_20;
  reg [31:0] _GEN_151;
  reg [9:0] accumulator_21;
  reg [31:0] _GEN_152;
  reg [9:0] accumulator_22;
  reg [31:0] _GEN_153;
  reg [9:0] accumulator_23;
  reg [31:0] _GEN_154;
  reg [9:0] accumulator_24;
  reg [31:0] _GEN_155;
  reg [9:0] accumulator_25;
  reg [31:0] _GEN_156;
  reg [9:0] accumulator_26;
  reg [31:0] _GEN_157;
  reg [9:0] accumulator_27;
  reg [31:0] _GEN_158;
  reg [9:0] accumulator_28;
  reg [31:0] _GEN_159;
  reg [9:0] accumulator_29;
  reg [31:0] _GEN_160;
  reg [9:0] accumulator_30;
  reg [31:0] _GEN_161;
  reg [9:0] accumulator_31;
  reg [31:0] _GEN_162;
  wire  _T_46;
  wire  _T_47;
  wire  _T_49;
  wire [9:0] _GEN_0;
  wire [9:0] _GEN_4;
  wire [9:0] _GEN_5;
  wire [9:0] _GEN_6;
  wire [9:0] _GEN_7;
  wire [9:0] _GEN_8;
  wire [9:0] _GEN_9;
  wire [9:0] _GEN_10;
  wire [9:0] _GEN_11;
  wire [9:0] _GEN_12;
  wire [9:0] _GEN_13;
  wire [9:0] _GEN_14;
  wire [9:0] _GEN_15;
  wire [9:0] _GEN_16;
  wire [9:0] _GEN_17;
  wire [9:0] _GEN_18;
  wire [9:0] _GEN_19;
  wire [9:0] _GEN_20;
  wire [9:0] _GEN_21;
  wire [9:0] _GEN_22;
  wire [9:0] _GEN_23;
  wire [9:0] _GEN_24;
  wire [9:0] _GEN_25;
  wire [9:0] _GEN_26;
  wire [9:0] _GEN_27;
  wire [9:0] _GEN_28;
  wire [9:0] _GEN_29;
  wire [9:0] _GEN_30;
  wire [9:0] _GEN_31;
  wire [9:0] _GEN_32;
  wire [9:0] _GEN_33;
  wire [9:0] _GEN_34;
  wire [9:0] _GEN_1;
  wire [10:0] _T_50;
  wire [9:0] _T_51;
  wire [9:0] _T_52;
  wire [9:0] _GEN_2;
  wire [9:0] _GEN_35;
  wire [9:0] _GEN_36;
  wire [9:0] _GEN_37;
  wire [9:0] _GEN_38;
  wire [9:0] _GEN_39;
  wire [9:0] _GEN_40;
  wire [9:0] _GEN_41;
  wire [9:0] _GEN_42;
  wire [9:0] _GEN_43;
  wire [9:0] _GEN_44;
  wire [9:0] _GEN_45;
  wire [9:0] _GEN_46;
  wire [9:0] _GEN_47;
  wire [9:0] _GEN_48;
  wire [9:0] _GEN_49;
  wire [9:0] _GEN_50;
  wire [9:0] _GEN_51;
  wire [9:0] _GEN_52;
  wire [9:0] _GEN_53;
  wire [9:0] _GEN_54;
  wire [9:0] _GEN_55;
  wire [9:0] _GEN_56;
  wire [9:0] _GEN_57;
  wire [9:0] _GEN_58;
  wire [9:0] _GEN_59;
  wire [9:0] _GEN_60;
  wire [9:0] _GEN_61;
  wire [9:0] _GEN_62;
  wire [9:0] _GEN_63;
  wire [9:0] _GEN_64;
  wire [9:0] _GEN_65;
  wire [9:0] _GEN_66;
  wire [9:0] _GEN_67;
  wire [9:0] _GEN_68;
  wire [9:0] _GEN_69;
  wire [9:0] _GEN_70;
  wire [9:0] _GEN_71;
  wire [9:0] _GEN_72;
  wire [9:0] _GEN_73;
  wire [9:0] _GEN_74;
  wire [9:0] _GEN_75;
  wire [9:0] _GEN_76;
  wire [9:0] _GEN_77;
  wire [9:0] _GEN_78;
  wire [9:0] _GEN_79;
  wire [9:0] _GEN_80;
  wire [9:0] _GEN_81;
  wire [9:0] _GEN_82;
  wire [9:0] _GEN_83;
  wire [9:0] _GEN_84;
  wire [9:0] _GEN_85;
  wire [9:0] _GEN_86;
  wire [9:0] _GEN_87;
  wire [9:0] _GEN_88;
  wire [9:0] _GEN_89;
  wire [9:0] _GEN_90;
  wire [9:0] _GEN_91;
  wire [9:0] _GEN_92;
  wire [9:0] _GEN_93;
  wire [9:0] _GEN_94;
  wire [9:0] _GEN_95;
  wire [9:0] _GEN_96;
  wire [9:0] _GEN_97;
  wire [9:0] _GEN_98;
  wire [9:0] _GEN_3;
  wire  _T_53;
  wire  _T_57;
  wire [9:0] _T_59;
  wire  _T_61;
  wire [9:0] _T_63;
  wire  _T_65;
  wire [9:0] _T_67;
  wire  _T_69;
  wire [9:0] _T_71;
  wire  _T_73;
  wire [9:0] _T_75;
  wire  _T_77;
  wire [9:0] _T_79;
  wire  _T_81;
  wire [9:0] _T_83;
  wire  _T_85;
  wire [9:0] _T_87;
  wire  _T_89;
  wire [9:0] _T_91;
  wire  _T_93;
  wire [9:0] _T_95;
  wire  _T_97;
  wire [9:0] _T_99;
  wire  _T_101;
  wire [9:0] _T_103;
  wire  _T_105;
  wire [9:0] _T_107;
  wire  _T_109;
  wire [9:0] _T_111;
  wire  _T_113;
  wire [9:0] _T_115;
  wire  _T_117;
  wire [9:0] _T_119;
  wire  _T_121;
  wire [9:0] _T_123;
  wire  _T_125;
  wire [9:0] _T_127;
  wire  _T_129;
  wire [9:0] _T_131;
  wire  _T_133;
  wire [9:0] _T_135;
  wire  _T_137;
  wire [9:0] _T_139;
  wire  _T_141;
  wire [9:0] _T_143;
  wire  _T_145;
  wire [9:0] _T_147;
  wire  _T_149;
  wire [9:0] _T_151;
  wire  _T_153;
  wire [9:0] _T_155;
  wire  _T_157;
  wire [9:0] _T_159;
  wire  _T_161;
  wire [9:0] _T_163;
  wire  _T_165;
  wire [9:0] _T_167;
  wire  _T_169;
  wire [9:0] _T_171;
  wire  _T_173;
  wire [9:0] _T_175;
  wire  _T_177;
  wire [9:0] _T_179;
  wire  _T_181;
  wire [9:0] _T_183;
  wire [9:0] _GEN_99;
  wire [9:0] _GEN_100;
  wire [9:0] _GEN_101;
  wire [9:0] _GEN_102;
  wire [9:0] _GEN_103;
  wire [9:0] _GEN_104;
  wire [9:0] _GEN_105;
  wire [9:0] _GEN_106;
  wire [9:0] _GEN_107;
  wire [9:0] _GEN_108;
  wire [9:0] _GEN_109;
  wire [9:0] _GEN_110;
  wire [9:0] _GEN_111;
  wire [9:0] _GEN_112;
  wire [9:0] _GEN_113;
  wire [9:0] _GEN_114;
  wire [9:0] _GEN_115;
  wire [9:0] _GEN_116;
  wire [9:0] _GEN_117;
  wire [9:0] _GEN_118;
  wire [9:0] _GEN_119;
  wire [9:0] _GEN_120;
  wire [9:0] _GEN_121;
  wire [9:0] _GEN_122;
  wire [9:0] _GEN_123;
  wire [9:0] _GEN_124;
  wire [9:0] _GEN_125;
  wire [9:0] _GEN_126;
  wire [9:0] _GEN_127;
  wire [9:0] _GEN_128;
  wire [9:0] _GEN_129;
  wire [9:0] _GEN_130;
  assign io_out = _GEN_3;
  assign _T_46 = io_reset == 1'h0;
  assign _T_47 = io_en & _T_46;
  assign _T_49 = reset == 1'h0;
  assign _GEN_0 = _GEN_34;
  assign _GEN_4 = 5'h1 == io_sel ? $signed(accumulator_1) : $signed(accumulator_0);
  assign _GEN_5 = 5'h2 == io_sel ? $signed(accumulator_2) : $signed(_GEN_4);
  assign _GEN_6 = 5'h3 == io_sel ? $signed(accumulator_3) : $signed(_GEN_5);
  assign _GEN_7 = 5'h4 == io_sel ? $signed(accumulator_4) : $signed(_GEN_6);
  assign _GEN_8 = 5'h5 == io_sel ? $signed(accumulator_5) : $signed(_GEN_7);
  assign _GEN_9 = 5'h6 == io_sel ? $signed(accumulator_6) : $signed(_GEN_8);
  assign _GEN_10 = 5'h7 == io_sel ? $signed(accumulator_7) : $signed(_GEN_9);
  assign _GEN_11 = 5'h8 == io_sel ? $signed(accumulator_8) : $signed(_GEN_10);
  assign _GEN_12 = 5'h9 == io_sel ? $signed(accumulator_9) : $signed(_GEN_11);
  assign _GEN_13 = 5'ha == io_sel ? $signed(accumulator_10) : $signed(_GEN_12);
  assign _GEN_14 = 5'hb == io_sel ? $signed(accumulator_11) : $signed(_GEN_13);
  assign _GEN_15 = 5'hc == io_sel ? $signed(accumulator_12) : $signed(_GEN_14);
  assign _GEN_16 = 5'hd == io_sel ? $signed(accumulator_13) : $signed(_GEN_15);
  assign _GEN_17 = 5'he == io_sel ? $signed(accumulator_14) : $signed(_GEN_16);
  assign _GEN_18 = 5'hf == io_sel ? $signed(accumulator_15) : $signed(_GEN_17);
  assign _GEN_19 = 5'h10 == io_sel ? $signed(accumulator_16) : $signed(_GEN_18);
  assign _GEN_20 = 5'h11 == io_sel ? $signed(accumulator_17) : $signed(_GEN_19);
  assign _GEN_21 = 5'h12 == io_sel ? $signed(accumulator_18) : $signed(_GEN_20);
  assign _GEN_22 = 5'h13 == io_sel ? $signed(accumulator_19) : $signed(_GEN_21);
  assign _GEN_23 = 5'h14 == io_sel ? $signed(accumulator_20) : $signed(_GEN_22);
  assign _GEN_24 = 5'h15 == io_sel ? $signed(accumulator_21) : $signed(_GEN_23);
  assign _GEN_25 = 5'h16 == io_sel ? $signed(accumulator_22) : $signed(_GEN_24);
  assign _GEN_26 = 5'h17 == io_sel ? $signed(accumulator_23) : $signed(_GEN_25);
  assign _GEN_27 = 5'h18 == io_sel ? $signed(accumulator_24) : $signed(_GEN_26);
  assign _GEN_28 = 5'h19 == io_sel ? $signed(accumulator_25) : $signed(_GEN_27);
  assign _GEN_29 = 5'h1a == io_sel ? $signed(accumulator_26) : $signed(_GEN_28);
  assign _GEN_30 = 5'h1b == io_sel ? $signed(accumulator_27) : $signed(_GEN_29);
  assign _GEN_31 = 5'h1c == io_sel ? $signed(accumulator_28) : $signed(_GEN_30);
  assign _GEN_32 = 5'h1d == io_sel ? $signed(accumulator_29) : $signed(_GEN_31);
  assign _GEN_33 = 5'h1e == io_sel ? $signed(accumulator_30) : $signed(_GEN_32);
  assign _GEN_34 = 5'h1f == io_sel ? $signed(accumulator_31) : $signed(_GEN_33);
  assign _GEN_1 = _GEN_34;
  assign _T_50 = $signed(_GEN_1) + $signed(io_in);
  assign _T_51 = _T_50[9:0];
  assign _T_52 = $signed(_T_51);
  assign _GEN_2 = _T_52;
  assign _GEN_35 = 5'h0 == io_sel ? $signed(_GEN_2) : $signed(accumulator_0);
  assign _GEN_36 = 5'h1 == io_sel ? $signed(_GEN_2) : $signed(accumulator_1);
  assign _GEN_37 = 5'h2 == io_sel ? $signed(_GEN_2) : $signed(accumulator_2);
  assign _GEN_38 = 5'h3 == io_sel ? $signed(_GEN_2) : $signed(accumulator_3);
  assign _GEN_39 = 5'h4 == io_sel ? $signed(_GEN_2) : $signed(accumulator_4);
  assign _GEN_40 = 5'h5 == io_sel ? $signed(_GEN_2) : $signed(accumulator_5);
  assign _GEN_41 = 5'h6 == io_sel ? $signed(_GEN_2) : $signed(accumulator_6);
  assign _GEN_42 = 5'h7 == io_sel ? $signed(_GEN_2) : $signed(accumulator_7);
  assign _GEN_43 = 5'h8 == io_sel ? $signed(_GEN_2) : $signed(accumulator_8);
  assign _GEN_44 = 5'h9 == io_sel ? $signed(_GEN_2) : $signed(accumulator_9);
  assign _GEN_45 = 5'ha == io_sel ? $signed(_GEN_2) : $signed(accumulator_10);
  assign _GEN_46 = 5'hb == io_sel ? $signed(_GEN_2) : $signed(accumulator_11);
  assign _GEN_47 = 5'hc == io_sel ? $signed(_GEN_2) : $signed(accumulator_12);
  assign _GEN_48 = 5'hd == io_sel ? $signed(_GEN_2) : $signed(accumulator_13);
  assign _GEN_49 = 5'he == io_sel ? $signed(_GEN_2) : $signed(accumulator_14);
  assign _GEN_50 = 5'hf == io_sel ? $signed(_GEN_2) : $signed(accumulator_15);
  assign _GEN_51 = 5'h10 == io_sel ? $signed(_GEN_2) : $signed(accumulator_16);
  assign _GEN_52 = 5'h11 == io_sel ? $signed(_GEN_2) : $signed(accumulator_17);
  assign _GEN_53 = 5'h12 == io_sel ? $signed(_GEN_2) : $signed(accumulator_18);
  assign _GEN_54 = 5'h13 == io_sel ? $signed(_GEN_2) : $signed(accumulator_19);
  assign _GEN_55 = 5'h14 == io_sel ? $signed(_GEN_2) : $signed(accumulator_20);
  assign _GEN_56 = 5'h15 == io_sel ? $signed(_GEN_2) : $signed(accumulator_21);
  assign _GEN_57 = 5'h16 == io_sel ? $signed(_GEN_2) : $signed(accumulator_22);
  assign _GEN_58 = 5'h17 == io_sel ? $signed(_GEN_2) : $signed(accumulator_23);
  assign _GEN_59 = 5'h18 == io_sel ? $signed(_GEN_2) : $signed(accumulator_24);
  assign _GEN_60 = 5'h19 == io_sel ? $signed(_GEN_2) : $signed(accumulator_25);
  assign _GEN_61 = 5'h1a == io_sel ? $signed(_GEN_2) : $signed(accumulator_26);
  assign _GEN_62 = 5'h1b == io_sel ? $signed(_GEN_2) : $signed(accumulator_27);
  assign _GEN_63 = 5'h1c == io_sel ? $signed(_GEN_2) : $signed(accumulator_28);
  assign _GEN_64 = 5'h1d == io_sel ? $signed(_GEN_2) : $signed(accumulator_29);
  assign _GEN_65 = 5'h1e == io_sel ? $signed(_GEN_2) : $signed(accumulator_30);
  assign _GEN_66 = 5'h1f == io_sel ? $signed(_GEN_2) : $signed(accumulator_31);
  assign _GEN_67 = _T_47 ? $signed(_GEN_35) : $signed(accumulator_0);
  assign _GEN_68 = _T_47 ? $signed(_GEN_36) : $signed(accumulator_1);
  assign _GEN_69 = _T_47 ? $signed(_GEN_37) : $signed(accumulator_2);
  assign _GEN_70 = _T_47 ? $signed(_GEN_38) : $signed(accumulator_3);
  assign _GEN_71 = _T_47 ? $signed(_GEN_39) : $signed(accumulator_4);
  assign _GEN_72 = _T_47 ? $signed(_GEN_40) : $signed(accumulator_5);
  assign _GEN_73 = _T_47 ? $signed(_GEN_41) : $signed(accumulator_6);
  assign _GEN_74 = _T_47 ? $signed(_GEN_42) : $signed(accumulator_7);
  assign _GEN_75 = _T_47 ? $signed(_GEN_43) : $signed(accumulator_8);
  assign _GEN_76 = _T_47 ? $signed(_GEN_44) : $signed(accumulator_9);
  assign _GEN_77 = _T_47 ? $signed(_GEN_45) : $signed(accumulator_10);
  assign _GEN_78 = _T_47 ? $signed(_GEN_46) : $signed(accumulator_11);
  assign _GEN_79 = _T_47 ? $signed(_GEN_47) : $signed(accumulator_12);
  assign _GEN_80 = _T_47 ? $signed(_GEN_48) : $signed(accumulator_13);
  assign _GEN_81 = _T_47 ? $signed(_GEN_49) : $signed(accumulator_14);
  assign _GEN_82 = _T_47 ? $signed(_GEN_50) : $signed(accumulator_15);
  assign _GEN_83 = _T_47 ? $signed(_GEN_51) : $signed(accumulator_16);
  assign _GEN_84 = _T_47 ? $signed(_GEN_52) : $signed(accumulator_17);
  assign _GEN_85 = _T_47 ? $signed(_GEN_53) : $signed(accumulator_18);
  assign _GEN_86 = _T_47 ? $signed(_GEN_54) : $signed(accumulator_19);
  assign _GEN_87 = _T_47 ? $signed(_GEN_55) : $signed(accumulator_20);
  assign _GEN_88 = _T_47 ? $signed(_GEN_56) : $signed(accumulator_21);
  assign _GEN_89 = _T_47 ? $signed(_GEN_57) : $signed(accumulator_22);
  assign _GEN_90 = _T_47 ? $signed(_GEN_58) : $signed(accumulator_23);
  assign _GEN_91 = _T_47 ? $signed(_GEN_59) : $signed(accumulator_24);
  assign _GEN_92 = _T_47 ? $signed(_GEN_60) : $signed(accumulator_25);
  assign _GEN_93 = _T_47 ? $signed(_GEN_61) : $signed(accumulator_26);
  assign _GEN_94 = _T_47 ? $signed(_GEN_62) : $signed(accumulator_27);
  assign _GEN_95 = _T_47 ? $signed(_GEN_63) : $signed(accumulator_28);
  assign _GEN_96 = _T_47 ? $signed(_GEN_64) : $signed(accumulator_29);
  assign _GEN_97 = _T_47 ? $signed(_GEN_65) : $signed(accumulator_30);
  assign _GEN_98 = _T_47 ? $signed(_GEN_66) : $signed(accumulator_31);
  assign _GEN_3 = _GEN_34;
  assign _T_53 = io_en & io_reset;
  assign _T_57 = 5'h0 == io_sel;
  assign _T_59 = _T_57 ? $signed(io_in) : $signed(10'sh0);
  assign _T_61 = 5'h1 == io_sel;
  assign _T_63 = _T_61 ? $signed(io_in) : $signed(10'sh0);
  assign _T_65 = 5'h2 == io_sel;
  assign _T_67 = _T_65 ? $signed(io_in) : $signed(10'sh0);
  assign _T_69 = 5'h3 == io_sel;
  assign _T_71 = _T_69 ? $signed(io_in) : $signed(10'sh0);
  assign _T_73 = 5'h4 == io_sel;
  assign _T_75 = _T_73 ? $signed(io_in) : $signed(10'sh0);
  assign _T_77 = 5'h5 == io_sel;
  assign _T_79 = _T_77 ? $signed(io_in) : $signed(10'sh0);
  assign _T_81 = 5'h6 == io_sel;
  assign _T_83 = _T_81 ? $signed(io_in) : $signed(10'sh0);
  assign _T_85 = 5'h7 == io_sel;
  assign _T_87 = _T_85 ? $signed(io_in) : $signed(10'sh0);
  assign _T_89 = 5'h8 == io_sel;
  assign _T_91 = _T_89 ? $signed(io_in) : $signed(10'sh0);
  assign _T_93 = 5'h9 == io_sel;
  assign _T_95 = _T_93 ? $signed(io_in) : $signed(10'sh0);
  assign _T_97 = 5'ha == io_sel;
  assign _T_99 = _T_97 ? $signed(io_in) : $signed(10'sh0);
  assign _T_101 = 5'hb == io_sel;
  assign _T_103 = _T_101 ? $signed(io_in) : $signed(10'sh0);
  assign _T_105 = 5'hc == io_sel;
  assign _T_107 = _T_105 ? $signed(io_in) : $signed(10'sh0);
  assign _T_109 = 5'hd == io_sel;
  assign _T_111 = _T_109 ? $signed(io_in) : $signed(10'sh0);
  assign _T_113 = 5'he == io_sel;
  assign _T_115 = _T_113 ? $signed(io_in) : $signed(10'sh0);
  assign _T_117 = 5'hf == io_sel;
  assign _T_119 = _T_117 ? $signed(io_in) : $signed(10'sh0);
  assign _T_121 = 5'h10 == io_sel;
  assign _T_123 = _T_121 ? $signed(io_in) : $signed(10'sh0);
  assign _T_125 = 5'h11 == io_sel;
  assign _T_127 = _T_125 ? $signed(io_in) : $signed(10'sh0);
  assign _T_129 = 5'h12 == io_sel;
  assign _T_131 = _T_129 ? $signed(io_in) : $signed(10'sh0);
  assign _T_133 = 5'h13 == io_sel;
  assign _T_135 = _T_133 ? $signed(io_in) : $signed(10'sh0);
  assign _T_137 = 5'h14 == io_sel;
  assign _T_139 = _T_137 ? $signed(io_in) : $signed(10'sh0);
  assign _T_141 = 5'h15 == io_sel;
  assign _T_143 = _T_141 ? $signed(io_in) : $signed(10'sh0);
  assign _T_145 = 5'h16 == io_sel;
  assign _T_147 = _T_145 ? $signed(io_in) : $signed(10'sh0);
  assign _T_149 = 5'h17 == io_sel;
  assign _T_151 = _T_149 ? $signed(io_in) : $signed(10'sh0);
  assign _T_153 = 5'h18 == io_sel;
  assign _T_155 = _T_153 ? $signed(io_in) : $signed(10'sh0);
  assign _T_157 = 5'h19 == io_sel;
  assign _T_159 = _T_157 ? $signed(io_in) : $signed(10'sh0);
  assign _T_161 = 5'h1a == io_sel;
  assign _T_163 = _T_161 ? $signed(io_in) : $signed(10'sh0);
  assign _T_165 = 5'h1b == io_sel;
  assign _T_167 = _T_165 ? $signed(io_in) : $signed(10'sh0);
  assign _T_169 = 5'h1c == io_sel;
  assign _T_171 = _T_169 ? $signed(io_in) : $signed(10'sh0);
  assign _T_173 = 5'h1d == io_sel;
  assign _T_175 = _T_173 ? $signed(io_in) : $signed(10'sh0);
  assign _T_177 = 5'h1e == io_sel;
  assign _T_179 = _T_177 ? $signed(io_in) : $signed(10'sh0);
  assign _T_181 = 5'h1f == io_sel;
  assign _T_183 = _T_181 ? $signed(io_in) : $signed(10'sh0);
  assign _GEN_99 = _T_53 ? $signed(_T_59) : $signed(_GEN_67);
  assign _GEN_100 = _T_53 ? $signed(_T_63) : $signed(_GEN_68);
  assign _GEN_101 = _T_53 ? $signed(_T_67) : $signed(_GEN_69);
  assign _GEN_102 = _T_53 ? $signed(_T_71) : $signed(_GEN_70);
  assign _GEN_103 = _T_53 ? $signed(_T_75) : $signed(_GEN_71);
  assign _GEN_104 = _T_53 ? $signed(_T_79) : $signed(_GEN_72);
  assign _GEN_105 = _T_53 ? $signed(_T_83) : $signed(_GEN_73);
  assign _GEN_106 = _T_53 ? $signed(_T_87) : $signed(_GEN_74);
  assign _GEN_107 = _T_53 ? $signed(_T_91) : $signed(_GEN_75);
  assign _GEN_108 = _T_53 ? $signed(_T_95) : $signed(_GEN_76);
  assign _GEN_109 = _T_53 ? $signed(_T_99) : $signed(_GEN_77);
  assign _GEN_110 = _T_53 ? $signed(_T_103) : $signed(_GEN_78);
  assign _GEN_111 = _T_53 ? $signed(_T_107) : $signed(_GEN_79);
  assign _GEN_112 = _T_53 ? $signed(_T_111) : $signed(_GEN_80);
  assign _GEN_113 = _T_53 ? $signed(_T_115) : $signed(_GEN_81);
  assign _GEN_114 = _T_53 ? $signed(_T_119) : $signed(_GEN_82);
  assign _GEN_115 = _T_53 ? $signed(_T_123) : $signed(_GEN_83);
  assign _GEN_116 = _T_53 ? $signed(_T_127) : $signed(_GEN_84);
  assign _GEN_117 = _T_53 ? $signed(_T_131) : $signed(_GEN_85);
  assign _GEN_118 = _T_53 ? $signed(_T_135) : $signed(_GEN_86);
  assign _GEN_119 = _T_53 ? $signed(_T_139) : $signed(_GEN_87);
  assign _GEN_120 = _T_53 ? $signed(_T_143) : $signed(_GEN_88);
  assign _GEN_121 = _T_53 ? $signed(_T_147) : $signed(_GEN_89);
  assign _GEN_122 = _T_53 ? $signed(_T_151) : $signed(_GEN_90);
  assign _GEN_123 = _T_53 ? $signed(_T_155) : $signed(_GEN_91);
  assign _GEN_124 = _T_53 ? $signed(_T_159) : $signed(_GEN_92);
  assign _GEN_125 = _T_53 ? $signed(_T_163) : $signed(_GEN_93);
  assign _GEN_126 = _T_53 ? $signed(_T_167) : $signed(_GEN_94);
  assign _GEN_127 = _T_53 ? $signed(_T_171) : $signed(_GEN_95);
  assign _GEN_128 = _T_53 ? $signed(_T_175) : $signed(_GEN_96);
  assign _GEN_129 = _T_53 ? $signed(_T_179) : $signed(_GEN_97);
  assign _GEN_130 = _T_53 ? $signed(_T_183) : $signed(_GEN_98);
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_131 = {1{$random}};
  accumulator_0 = _GEN_131[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_132 = {1{$random}};
  accumulator_1 = _GEN_132[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_133 = {1{$random}};
  accumulator_2 = _GEN_133[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_134 = {1{$random}};
  accumulator_3 = _GEN_134[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_135 = {1{$random}};
  accumulator_4 = _GEN_135[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_136 = {1{$random}};
  accumulator_5 = _GEN_136[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_137 = {1{$random}};
  accumulator_6 = _GEN_137[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_138 = {1{$random}};
  accumulator_7 = _GEN_138[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_139 = {1{$random}};
  accumulator_8 = _GEN_139[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_140 = {1{$random}};
  accumulator_9 = _GEN_140[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_141 = {1{$random}};
  accumulator_10 = _GEN_141[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_142 = {1{$random}};
  accumulator_11 = _GEN_142[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_143 = {1{$random}};
  accumulator_12 = _GEN_143[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_144 = {1{$random}};
  accumulator_13 = _GEN_144[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_145 = {1{$random}};
  accumulator_14 = _GEN_145[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_146 = {1{$random}};
  accumulator_15 = _GEN_146[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_147 = {1{$random}};
  accumulator_16 = _GEN_147[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_148 = {1{$random}};
  accumulator_17 = _GEN_148[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_149 = {1{$random}};
  accumulator_18 = _GEN_149[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_150 = {1{$random}};
  accumulator_19 = _GEN_150[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_151 = {1{$random}};
  accumulator_20 = _GEN_151[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_152 = {1{$random}};
  accumulator_21 = _GEN_152[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_153 = {1{$random}};
  accumulator_22 = _GEN_153[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_154 = {1{$random}};
  accumulator_23 = _GEN_154[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_155 = {1{$random}};
  accumulator_24 = _GEN_155[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_156 = {1{$random}};
  accumulator_25 = _GEN_156[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_157 = {1{$random}};
  accumulator_26 = _GEN_157[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_158 = {1{$random}};
  accumulator_27 = _GEN_158[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_159 = {1{$random}};
  accumulator_28 = _GEN_159[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_160 = {1{$random}};
  accumulator_29 = _GEN_160[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_161 = {1{$random}};
  accumulator_30 = _GEN_161[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_162 = {1{$random}};
  accumulator_31 = _GEN_162[9:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (_T_53) begin
      if (_T_57) begin
        accumulator_0 <= io_in;
      end else begin
        accumulator_0 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h0 == io_sel) begin
          accumulator_0 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_61) begin
        accumulator_1 <= io_in;
      end else begin
        accumulator_1 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h1 == io_sel) begin
          accumulator_1 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_65) begin
        accumulator_2 <= io_in;
      end else begin
        accumulator_2 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h2 == io_sel) begin
          accumulator_2 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_69) begin
        accumulator_3 <= io_in;
      end else begin
        accumulator_3 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h3 == io_sel) begin
          accumulator_3 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_73) begin
        accumulator_4 <= io_in;
      end else begin
        accumulator_4 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h4 == io_sel) begin
          accumulator_4 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_77) begin
        accumulator_5 <= io_in;
      end else begin
        accumulator_5 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h5 == io_sel) begin
          accumulator_5 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_81) begin
        accumulator_6 <= io_in;
      end else begin
        accumulator_6 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h6 == io_sel) begin
          accumulator_6 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_85) begin
        accumulator_7 <= io_in;
      end else begin
        accumulator_7 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h7 == io_sel) begin
          accumulator_7 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_89) begin
        accumulator_8 <= io_in;
      end else begin
        accumulator_8 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h8 == io_sel) begin
          accumulator_8 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_93) begin
        accumulator_9 <= io_in;
      end else begin
        accumulator_9 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h9 == io_sel) begin
          accumulator_9 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_97) begin
        accumulator_10 <= io_in;
      end else begin
        accumulator_10 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'ha == io_sel) begin
          accumulator_10 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_101) begin
        accumulator_11 <= io_in;
      end else begin
        accumulator_11 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'hb == io_sel) begin
          accumulator_11 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_105) begin
        accumulator_12 <= io_in;
      end else begin
        accumulator_12 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'hc == io_sel) begin
          accumulator_12 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_109) begin
        accumulator_13 <= io_in;
      end else begin
        accumulator_13 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'hd == io_sel) begin
          accumulator_13 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_113) begin
        accumulator_14 <= io_in;
      end else begin
        accumulator_14 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'he == io_sel) begin
          accumulator_14 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_117) begin
        accumulator_15 <= io_in;
      end else begin
        accumulator_15 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'hf == io_sel) begin
          accumulator_15 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_121) begin
        accumulator_16 <= io_in;
      end else begin
        accumulator_16 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h10 == io_sel) begin
          accumulator_16 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_125) begin
        accumulator_17 <= io_in;
      end else begin
        accumulator_17 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h11 == io_sel) begin
          accumulator_17 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_129) begin
        accumulator_18 <= io_in;
      end else begin
        accumulator_18 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h12 == io_sel) begin
          accumulator_18 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_133) begin
        accumulator_19 <= io_in;
      end else begin
        accumulator_19 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h13 == io_sel) begin
          accumulator_19 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_137) begin
        accumulator_20 <= io_in;
      end else begin
        accumulator_20 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h14 == io_sel) begin
          accumulator_20 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_141) begin
        accumulator_21 <= io_in;
      end else begin
        accumulator_21 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h15 == io_sel) begin
          accumulator_21 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_145) begin
        accumulator_22 <= io_in;
      end else begin
        accumulator_22 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h16 == io_sel) begin
          accumulator_22 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_149) begin
        accumulator_23 <= io_in;
      end else begin
        accumulator_23 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h17 == io_sel) begin
          accumulator_23 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_153) begin
        accumulator_24 <= io_in;
      end else begin
        accumulator_24 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h18 == io_sel) begin
          accumulator_24 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_157) begin
        accumulator_25 <= io_in;
      end else begin
        accumulator_25 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h19 == io_sel) begin
          accumulator_25 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_161) begin
        accumulator_26 <= io_in;
      end else begin
        accumulator_26 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h1a == io_sel) begin
          accumulator_26 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_165) begin
        accumulator_27 <= io_in;
      end else begin
        accumulator_27 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h1b == io_sel) begin
          accumulator_27 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_169) begin
        accumulator_28 <= io_in;
      end else begin
        accumulator_28 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h1c == io_sel) begin
          accumulator_28 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_173) begin
        accumulator_29 <= io_in;
      end else begin
        accumulator_29 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h1d == io_sel) begin
          accumulator_29 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_177) begin
        accumulator_30 <= io_in;
      end else begin
        accumulator_30 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h1e == io_sel) begin
          accumulator_30 <= _GEN_2;
        end
      end
    end
    if (_T_53) begin
      if (_T_181) begin
        accumulator_31 <= io_in;
      end else begin
        accumulator_31 <= 10'sh0;
      end
    end else begin
      if (_T_47) begin
        if (5'h1f == io_sel) begin
          accumulator_31 <= _GEN_2;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_47 & _T_49) begin
          $fwrite(32'h80000002,"Acc Update! %d, %d, %d\n",io_in,_GEN_0,io_sel);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_49) begin
          $fwrite(32'h80000002,"Acc Reset! %d @ %d\n",io_in,io_sel);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module MulAdd(
  input  [15:0] io_a,
  input  [9:0]  io_b,
  input  [31:0] io_m,
  input  [15:0] io_c,
  output [31:0] io_r
);
  wire [15:0] _GEN_0;
  wire [25:0] _T_7;
  wire [32:0] _T_8;
  wire [32:0] _GEN_1;
  wire [58:0] _T_9;
  wire [57:0] _T_10;
  wire [57:0] _T_11;
  wire [57:0] _GEN_2;
  wire [58:0] _T_12;
  wire [57:0] _T_13;
  wire [57:0] _T_14;
  wire [31:0] _GEN_3;
  assign io_r = $signed(_GEN_3);
  assign _GEN_0 = {{6{io_b[9]}},io_b};
  assign _T_7 = $signed(io_a) * $signed(_GEN_0);
  assign _T_8 = {1'b0,$signed(io_m)};
  assign _GEN_1 = {{7{_T_7[25]}},_T_7};
  assign _T_9 = $signed(_GEN_1) * $signed(_T_8);
  assign _T_10 = _T_9[57:0];
  assign _T_11 = $signed(_T_10);
  assign _GEN_2 = {{42{io_c[15]}},io_c};
  assign _T_12 = $signed(_T_11) + $signed(_GEN_2);
  assign _T_13 = _T_12[57:0];
  assign _T_14 = $signed(_T_13);
  assign _GEN_3 = _T_14[31:0];
endmodule
module XNORNetInference(
  input          clock,
  input          reset,
  input  [127:0] io_input,
  input          io_inputPush,
  input          io_inputBufferPush,
  input          io_inputBufferPop,
  input          io_inputBufferReset,
  input  [7:0]   io_memAddr,
  output [127:0] io_memOut,
  input          io_memWen,
  input  [127:0] io_memIn,
  input  [7:0]   io_memWAddr,
  input          io_accEn,
  input  [4:0]   io_accSel,
  input          io_accReset,
  input          io_maxReset,
  input          io_maxEn,
  input  [3:0]   io_maxOffset,
  input  [15:0]  io_featureNumInverse65536,
  input  [15:0]  io_actualFeatureNum,
  input          io_meanReset,
  input          io_meanUpdate,
  input          io_meanBufferReset,
  output [3:0]   io_result,
  output [31:0]  io_mean,
  output [15:0]  io_maa,
  output [15:0]  io_mab,
  output [31:0]  io_mam,
  output [15:0]  io_mac
);
  wire  mem_clock;
  wire [7:0] mem_io_addr;
  wire [7:0] mem_io_waddr;
  wire [127:0] mem_io_in;
  wire [127:0] mem_io_out;
  wire  mem_io_wen;
  wire  mem_io_ren;
  wire [3:0] inputWire;
  wire  binaryBuffer_clock;
  wire  binaryBuffer_io_reset;
  wire [3:0] binaryBuffer_io_in;
  wire [127:0] binaryBuffer_io_fastin;
  wire  binaryBuffer_io_push;
  wire  binaryBuffer_io_fastpush;
  wire [31:0] binaryBuffer_io_out;
  wire  binaryBuffer_io_pop;
  wire [31:0] xnor$_io_in1;
  wire [31:0] xnor$_io_in2_0;
  wire [31:0] xnor$_io_in2_1;
  wire [31:0] xnor$_io_in2_2;
  wire [31:0] xnor$_io_in2_3;
  wire [31:0] xnor$_io_out_0;
  wire [31:0] xnor$_io_out_1;
  wire [31:0] xnor$_io_out_2;
  wire [31:0] xnor$_io_out_3;
  wire [127:0] _T_33;
  wire [31:0] _T_44_0;
  wire [31:0] _T_44_1;
  wire [31:0] _T_44_2;
  wire [31:0] _T_44_3;
  wire [127:0] _T_57;
  wire [31:0] _T_58;
  wire [31:0] _T_59;
  wire [31:0] _T_60;
  wire [31:0] _T_61;
  wire  meanBuffer_clock;
  wire [31:0] meanBuffer_io_in_0;
  wire [31:0] meanBuffer_io_in_1;
  wire [31:0] meanBuffer_io_in_2;
  wire [31:0] meanBuffer_io_in_3;
  wire [15:0] meanBuffer_io_cntInverse65536;
  wire  meanBuffer_io_reset;
  wire [31:0] meanBuffer_io_out;
  wire  mean_clock;
  wire  mean_reset;
  wire  mean_io_reset;
  wire [31:0] mean_io_input;
  wire  mean_io_update;
  wire [31:0] mean_io_output;
  wire  maxModule_clock;
  wire  maxModule_io_reset;
  wire  maxModule_io_en;
  wire [31:0] maxModule_io_in_0;
  wire [31:0] maxModule_io_in_1;
  wire [31:0] maxModule_io_in_2;
  wire [31:0] maxModule_io_in_3;
  wire [3:0] maxModule_io_offset;
  wire [3:0] maxModule_io_out;
  wire [3:0] maxModule_io_maxLen;
  wire  Accumulator_clock;
  wire  Accumulator_reset;
  wire [9:0] Accumulator_io_in;
  wire [9:0] Accumulator_io_out;
  wire [4:0] Accumulator_io_sel;
  wire  Accumulator_io_en;
  wire  Accumulator_io_reset;
  wire [3:0] _T_62;
  wire [3:0] _T_63;
  wire [3:0] _T_64;
  wire [3:0] _T_65;
  wire [3:0] _T_66;
  wire [3:0] _T_67;
  wire [3:0] _T_68;
  wire [3:0] _T_69;
  reg [5:0] _T_72;
  reg [31:0] _GEN_518;
  reg [5:0] _T_75;
  reg [31:0] _GEN_519;
  reg [5:0] _T_78;
  reg [31:0] _GEN_520;
  reg [5:0] _T_81;
  reg [31:0] _GEN_521;
  reg [5:0] _T_84;
  reg [31:0] _GEN_522;
  reg [5:0] _T_87;
  reg [31:0] _GEN_523;
  reg [5:0] _T_90;
  reg [31:0] _GEN_524;
  reg [5:0] _T_93;
  reg [31:0] _GEN_525;
  reg [5:0] _T_96;
  reg [31:0] _GEN_526;
  reg [5:0] _T_99;
  reg [31:0] _GEN_527;
  reg [5:0] _T_102;
  reg [31:0] _GEN_528;
  reg [5:0] _T_105;
  reg [31:0] _GEN_529;
  reg [5:0] _T_108;
  reg [31:0] _GEN_530;
  reg [5:0] _T_111;
  reg [31:0] _GEN_531;
  reg [5:0] _T_114;
  reg [31:0] _GEN_532;
  reg [5:0] _T_117;
  reg [31:0] _GEN_533;
  wire [5:0] _T_120_0;
  wire [5:0] _T_120_1;
  wire [5:0] _T_120_2;
  wire [5:0] _T_120_3;
  wire [5:0] _T_120_4;
  wire [5:0] _T_120_5;
  wire [5:0] _T_120_6;
  wire [5:0] _T_120_7;
  wire [5:0] _T_120_8;
  wire [5:0] _T_120_9;
  wire [5:0] _T_120_10;
  wire [5:0] _T_120_11;
  wire [5:0] _T_120_12;
  wire [5:0] _T_120_13;
  wire [5:0] _T_120_14;
  wire [5:0] _T_120_15;
  reg [5:0] _T_142;
  reg [31:0] _GEN_534;
  reg [5:0] _T_145;
  reg [31:0] _GEN_535;
  reg [5:0] _T_148;
  reg [31:0] _GEN_536;
  reg [5:0] _T_151;
  reg [31:0] _GEN_537;
  reg [5:0] _T_154;
  reg [31:0] _GEN_538;
  reg [5:0] _T_157;
  reg [31:0] _GEN_539;
  reg [5:0] _T_160;
  reg [31:0] _GEN_540;
  reg [5:0] _T_163;
  reg [31:0] _GEN_541;
  reg [5:0] _T_166;
  reg [31:0] _GEN_542;
  reg [5:0] _T_169;
  reg [31:0] _GEN_543;
  reg [5:0] _T_172;
  reg [31:0] _GEN_544;
  reg [5:0] _T_175;
  reg [31:0] _GEN_545;
  reg [5:0] _T_178;
  reg [31:0] _GEN_546;
  reg [5:0] _T_181;
  reg [31:0] _GEN_547;
  reg [5:0] _T_184;
  reg [31:0] _GEN_548;
  reg [5:0] _T_187;
  reg [31:0] _GEN_549;
  wire [5:0] _T_190_0;
  wire [5:0] _T_190_1;
  wire [5:0] _T_190_2;
  wire [5:0] _T_190_3;
  wire [5:0] _T_190_4;
  wire [5:0] _T_190_5;
  wire [5:0] _T_190_6;
  wire [5:0] _T_190_7;
  wire [5:0] _T_190_8;
  wire [5:0] _T_190_9;
  wire [5:0] _T_190_10;
  wire [5:0] _T_190_11;
  wire [5:0] _T_190_12;
  wire [5:0] _T_190_13;
  wire [5:0] _T_190_14;
  wire [5:0] _T_190_15;
  reg [5:0] _T_212;
  reg [31:0] _GEN_550;
  reg [5:0] _T_215;
  reg [31:0] _GEN_551;
  reg [5:0] _T_218;
  reg [31:0] _GEN_552;
  reg [5:0] _T_221;
  reg [31:0] _GEN_553;
  reg [5:0] _T_224;
  reg [31:0] _GEN_554;
  reg [5:0] _T_227;
  reg [31:0] _GEN_555;
  reg [5:0] _T_230;
  reg [31:0] _GEN_556;
  reg [5:0] _T_233;
  reg [31:0] _GEN_557;
  reg [5:0] _T_236;
  reg [31:0] _GEN_558;
  reg [5:0] _T_239;
  reg [31:0] _GEN_559;
  reg [5:0] _T_242;
  reg [31:0] _GEN_560;
  reg [5:0] _T_245;
  reg [31:0] _GEN_561;
  reg [5:0] _T_248;
  reg [31:0] _GEN_562;
  reg [5:0] _T_251;
  reg [31:0] _GEN_563;
  reg [5:0] _T_254;
  reg [31:0] _GEN_564;
  reg [5:0] _T_257;
  reg [31:0] _GEN_565;
  wire [5:0] _T_260_0;
  wire [5:0] _T_260_1;
  wire [5:0] _T_260_2;
  wire [5:0] _T_260_3;
  wire [5:0] _T_260_4;
  wire [5:0] _T_260_5;
  wire [5:0] _T_260_6;
  wire [5:0] _T_260_7;
  wire [5:0] _T_260_8;
  wire [5:0] _T_260_9;
  wire [5:0] _T_260_10;
  wire [5:0] _T_260_11;
  wire [5:0] _T_260_12;
  wire [5:0] _T_260_13;
  wire [5:0] _T_260_14;
  wire [5:0] _T_260_15;
  reg [5:0] _T_282;
  reg [31:0] _GEN_566;
  reg [5:0] _T_285;
  reg [31:0] _GEN_567;
  reg [5:0] _T_288;
  reg [31:0] _GEN_568;
  reg [5:0] _T_291;
  reg [31:0] _GEN_569;
  reg [5:0] _T_294;
  reg [31:0] _GEN_570;
  reg [5:0] _T_297;
  reg [31:0] _GEN_571;
  reg [5:0] _T_300;
  reg [31:0] _GEN_572;
  reg [5:0] _T_303;
  reg [31:0] _GEN_573;
  reg [5:0] _T_306;
  reg [31:0] _GEN_574;
  reg [5:0] _T_309;
  reg [31:0] _GEN_575;
  reg [5:0] _T_312;
  reg [31:0] _GEN_576;
  reg [5:0] _T_315;
  reg [31:0] _GEN_577;
  reg [5:0] _T_318;
  reg [31:0] _GEN_578;
  reg [5:0] _T_321;
  reg [31:0] _GEN_579;
  reg [5:0] _T_324;
  reg [31:0] _GEN_580;
  reg [5:0] _T_327;
  reg [31:0] _GEN_581;
  wire [5:0] _T_330_0;
  wire [5:0] _T_330_1;
  wire [5:0] _T_330_2;
  wire [5:0] _T_330_3;
  wire [5:0] _T_330_4;
  wire [5:0] _T_330_5;
  wire [5:0] _T_330_6;
  wire [5:0] _T_330_7;
  wire [5:0] _T_330_8;
  wire [5:0] _T_330_9;
  wire [5:0] _T_330_10;
  wire [5:0] _T_330_11;
  wire [5:0] _T_330_12;
  wire [5:0] _T_330_13;
  wire [5:0] _T_330_14;
  wire [5:0] _T_330_15;
  reg [5:0] _T_352;
  reg [31:0] _GEN_582;
  reg [5:0] _T_355;
  reg [31:0] _GEN_583;
  reg [5:0] _T_358;
  reg [31:0] _GEN_584;
  reg [5:0] _T_361;
  reg [31:0] _GEN_585;
  reg [5:0] _T_364;
  reg [31:0] _GEN_586;
  reg [5:0] _T_367;
  reg [31:0] _GEN_587;
  reg [5:0] _T_370;
  reg [31:0] _GEN_588;
  reg [5:0] _T_373;
  reg [31:0] _GEN_589;
  reg [5:0] _T_376;
  reg [31:0] _GEN_590;
  reg [5:0] _T_379;
  reg [31:0] _GEN_591;
  reg [5:0] _T_382;
  reg [31:0] _GEN_592;
  reg [5:0] _T_385;
  reg [31:0] _GEN_593;
  reg [5:0] _T_388;
  reg [31:0] _GEN_594;
  reg [5:0] _T_391;
  reg [31:0] _GEN_595;
  reg [5:0] _T_394;
  reg [31:0] _GEN_596;
  reg [5:0] _T_397;
  reg [31:0] _GEN_597;
  wire [5:0] _T_400_0;
  wire [5:0] _T_400_1;
  wire [5:0] _T_400_2;
  wire [5:0] _T_400_3;
  wire [5:0] _T_400_4;
  wire [5:0] _T_400_5;
  wire [5:0] _T_400_6;
  wire [5:0] _T_400_7;
  wire [5:0] _T_400_8;
  wire [5:0] _T_400_9;
  wire [5:0] _T_400_10;
  wire [5:0] _T_400_11;
  wire [5:0] _T_400_12;
  wire [5:0] _T_400_13;
  wire [5:0] _T_400_14;
  wire [5:0] _T_400_15;
  reg [5:0] _T_422;
  reg [31:0] _GEN_598;
  reg [5:0] _T_425;
  reg [31:0] _GEN_599;
  reg [5:0] _T_428;
  reg [31:0] _GEN_600;
  reg [5:0] _T_431;
  reg [31:0] _GEN_601;
  reg [5:0] _T_434;
  reg [31:0] _GEN_602;
  reg [5:0] _T_437;
  reg [31:0] _GEN_603;
  reg [5:0] _T_440;
  reg [31:0] _GEN_604;
  reg [5:0] _T_443;
  reg [31:0] _GEN_605;
  reg [5:0] _T_446;
  reg [31:0] _GEN_606;
  reg [5:0] _T_449;
  reg [31:0] _GEN_607;
  reg [5:0] _T_452;
  reg [31:0] _GEN_608;
  reg [5:0] _T_455;
  reg [31:0] _GEN_609;
  reg [5:0] _T_458;
  reg [31:0] _GEN_610;
  reg [5:0] _T_461;
  reg [31:0] _GEN_611;
  reg [5:0] _T_464;
  reg [31:0] _GEN_612;
  reg [5:0] _T_467;
  reg [31:0] _GEN_613;
  wire [5:0] _T_470_0;
  wire [5:0] _T_470_1;
  wire [5:0] _T_470_2;
  wire [5:0] _T_470_3;
  wire [5:0] _T_470_4;
  wire [5:0] _T_470_5;
  wire [5:0] _T_470_6;
  wire [5:0] _T_470_7;
  wire [5:0] _T_470_8;
  wire [5:0] _T_470_9;
  wire [5:0] _T_470_10;
  wire [5:0] _T_470_11;
  wire [5:0] _T_470_12;
  wire [5:0] _T_470_13;
  wire [5:0] _T_470_14;
  wire [5:0] _T_470_15;
  reg [5:0] _T_492;
  reg [31:0] _GEN_614;
  reg [5:0] _T_495;
  reg [31:0] _GEN_615;
  reg [5:0] _T_498;
  reg [31:0] _GEN_616;
  reg [5:0] _T_501;
  reg [31:0] _GEN_617;
  reg [5:0] _T_504;
  reg [31:0] _GEN_618;
  reg [5:0] _T_507;
  reg [31:0] _GEN_619;
  reg [5:0] _T_510;
  reg [31:0] _GEN_620;
  reg [5:0] _T_513;
  reg [31:0] _GEN_621;
  reg [5:0] _T_516;
  reg [31:0] _GEN_622;
  reg [5:0] _T_519;
  reg [31:0] _GEN_623;
  reg [5:0] _T_522;
  reg [31:0] _GEN_624;
  reg [5:0] _T_525;
  reg [31:0] _GEN_625;
  reg [5:0] _T_528;
  reg [31:0] _GEN_626;
  reg [5:0] _T_531;
  reg [31:0] _GEN_627;
  reg [5:0] _T_534;
  reg [31:0] _GEN_628;
  reg [5:0] _T_537;
  reg [31:0] _GEN_629;
  wire [5:0] _T_540_0;
  wire [5:0] _T_540_1;
  wire [5:0] _T_540_2;
  wire [5:0] _T_540_3;
  wire [5:0] _T_540_4;
  wire [5:0] _T_540_5;
  wire [5:0] _T_540_6;
  wire [5:0] _T_540_7;
  wire [5:0] _T_540_8;
  wire [5:0] _T_540_9;
  wire [5:0] _T_540_10;
  wire [5:0] _T_540_11;
  wire [5:0] _T_540_12;
  wire [5:0] _T_540_13;
  wire [5:0] _T_540_14;
  wire [5:0] _T_540_15;
  reg [5:0] _T_562;
  reg [31:0] _GEN_630;
  reg [5:0] _T_565;
  reg [31:0] _GEN_631;
  reg [5:0] _T_568;
  reg [31:0] _GEN_632;
  reg [5:0] _T_571;
  reg [31:0] _GEN_633;
  reg [5:0] _T_574;
  reg [31:0] _GEN_634;
  reg [5:0] _T_577;
  reg [31:0] _GEN_635;
  reg [5:0] _T_580;
  reg [31:0] _GEN_636;
  reg [5:0] _T_583;
  reg [31:0] _GEN_637;
  reg [5:0] _T_586;
  reg [31:0] _GEN_638;
  reg [5:0] _T_589;
  reg [31:0] _GEN_639;
  reg [5:0] _T_592;
  reg [31:0] _GEN_640;
  reg [5:0] _T_595;
  reg [31:0] _GEN_641;
  reg [5:0] _T_598;
  reg [31:0] _GEN_642;
  reg [5:0] _T_601;
  reg [31:0] _GEN_643;
  reg [5:0] _T_604;
  reg [31:0] _GEN_644;
  reg [5:0] _T_607;
  reg [31:0] _GEN_645;
  wire [5:0] _T_610_0;
  wire [5:0] _T_610_1;
  wire [5:0] _T_610_2;
  wire [5:0] _T_610_3;
  wire [5:0] _T_610_4;
  wire [5:0] _T_610_5;
  wire [5:0] _T_610_6;
  wire [5:0] _T_610_7;
  wire [5:0] _T_610_8;
  wire [5:0] _T_610_9;
  wire [5:0] _T_610_10;
  wire [5:0] _T_610_11;
  wire [5:0] _T_610_12;
  wire [5:0] _T_610_13;
  wire [5:0] _T_610_14;
  wire [5:0] _T_610_15;
  wire [5:0] _GEN_0;
  wire [5:0] _GEN_32;
  wire [5:0] _GEN_33;
  wire [5:0] _GEN_34;
  wire [5:0] _GEN_35;
  wire [5:0] _GEN_36;
  wire [5:0] _GEN_37;
  wire [5:0] _GEN_38;
  wire [5:0] _GEN_39;
  wire [5:0] _GEN_40;
  wire [5:0] _GEN_41;
  wire [5:0] _GEN_42;
  wire [5:0] _GEN_43;
  wire [5:0] _GEN_44;
  wire [5:0] _GEN_45;
  wire [5:0] _GEN_46;
  wire [5:0] _GEN_1;
  wire [5:0] _GEN_47;
  wire [5:0] _GEN_48;
  wire [5:0] _GEN_49;
  wire [5:0] _GEN_50;
  wire [5:0] _GEN_51;
  wire [5:0] _GEN_52;
  wire [5:0] _GEN_53;
  wire [5:0] _GEN_54;
  wire [5:0] _GEN_55;
  wire [5:0] _GEN_56;
  wire [5:0] _GEN_57;
  wire [5:0] _GEN_58;
  wire [5:0] _GEN_59;
  wire [5:0] _GEN_60;
  wire [5:0] _GEN_61;
  wire [6:0] _T_630;
  wire [5:0] _T_631;
  wire [5:0] _T_632;
  wire [5:0] _GEN_2;
  wire [5:0] _GEN_62;
  wire [5:0] _GEN_63;
  wire [5:0] _GEN_64;
  wire [5:0] _GEN_65;
  wire [5:0] _GEN_66;
  wire [5:0] _GEN_67;
  wire [5:0] _GEN_68;
  wire [5:0] _GEN_69;
  wire [5:0] _GEN_70;
  wire [5:0] _GEN_71;
  wire [5:0] _GEN_72;
  wire [5:0] _GEN_73;
  wire [5:0] _GEN_74;
  wire [5:0] _GEN_75;
  wire [5:0] _GEN_76;
  wire [5:0] _GEN_3;
  wire [5:0] _GEN_77;
  wire [5:0] _GEN_78;
  wire [5:0] _GEN_79;
  wire [5:0] _GEN_80;
  wire [5:0] _GEN_81;
  wire [5:0] _GEN_82;
  wire [5:0] _GEN_83;
  wire [5:0] _GEN_84;
  wire [5:0] _GEN_85;
  wire [5:0] _GEN_86;
  wire [5:0] _GEN_87;
  wire [5:0] _GEN_88;
  wire [5:0] _GEN_89;
  wire [5:0] _GEN_90;
  wire [5:0] _GEN_91;
  wire [6:0] _T_633;
  wire [5:0] _T_634;
  wire [5:0] _T_635;
  wire [5:0] _GEN_4;
  wire [5:0] _GEN_92;
  wire [5:0] _GEN_93;
  wire [5:0] _GEN_94;
  wire [5:0] _GEN_95;
  wire [5:0] _GEN_96;
  wire [5:0] _GEN_97;
  wire [5:0] _GEN_98;
  wire [5:0] _GEN_99;
  wire [5:0] _GEN_100;
  wire [5:0] _GEN_101;
  wire [5:0] _GEN_102;
  wire [5:0] _GEN_103;
  wire [5:0] _GEN_104;
  wire [5:0] _GEN_105;
  wire [5:0] _GEN_106;
  wire [5:0] _GEN_5;
  wire [5:0] _GEN_107;
  wire [5:0] _GEN_108;
  wire [5:0] _GEN_109;
  wire [5:0] _GEN_110;
  wire [5:0] _GEN_111;
  wire [5:0] _GEN_112;
  wire [5:0] _GEN_113;
  wire [5:0] _GEN_114;
  wire [5:0] _GEN_115;
  wire [5:0] _GEN_116;
  wire [5:0] _GEN_117;
  wire [5:0] _GEN_118;
  wire [5:0] _GEN_119;
  wire [5:0] _GEN_120;
  wire [5:0] _GEN_121;
  wire [6:0] _T_636;
  wire [5:0] _T_637;
  wire [5:0] _T_638;
  wire [5:0] _GEN_6;
  wire [5:0] _GEN_122;
  wire [5:0] _GEN_123;
  wire [5:0] _GEN_124;
  wire [5:0] _GEN_125;
  wire [5:0] _GEN_126;
  wire [5:0] _GEN_127;
  wire [5:0] _GEN_128;
  wire [5:0] _GEN_129;
  wire [5:0] _GEN_130;
  wire [5:0] _GEN_131;
  wire [5:0] _GEN_132;
  wire [5:0] _GEN_133;
  wire [5:0] _GEN_134;
  wire [5:0] _GEN_135;
  wire [5:0] _GEN_136;
  wire [5:0] _GEN_7;
  wire [5:0] _GEN_137;
  wire [5:0] _GEN_138;
  wire [5:0] _GEN_139;
  wire [5:0] _GEN_140;
  wire [5:0] _GEN_141;
  wire [5:0] _GEN_142;
  wire [5:0] _GEN_143;
  wire [5:0] _GEN_144;
  wire [5:0] _GEN_145;
  wire [5:0] _GEN_146;
  wire [5:0] _GEN_147;
  wire [5:0] _GEN_148;
  wire [5:0] _GEN_149;
  wire [5:0] _GEN_150;
  wire [5:0] _GEN_151;
  wire [6:0] _T_639;
  wire [5:0] _T_640;
  wire [5:0] _T_641;
  wire [6:0] _T_642;
  wire [5:0] _T_643;
  wire [5:0] _T_644;
  wire [6:0] _T_645;
  wire [5:0] _T_646;
  wire [5:0] _T_647;
  wire [6:0] _T_648;
  wire [5:0] _T_649;
  wire [5:0] _T_650;
  wire [15:0] MulAdd_io_a;
  wire [9:0] MulAdd_io_b;
  wire [31:0] MulAdd_io_m;
  wire [15:0] MulAdd_io_c;
  wire [31:0] MulAdd_io_r;
  wire [31:0] _T_651;
  wire [15:0] _T_652;
  wire [15:0] _T_653;
  wire [15:0] _T_654;
  wire [15:0] _T_655;
  wire  _T_656;
  wire  signs_0;
  wire  Accumulator_1_clock;
  wire  Accumulator_1_reset;
  wire [9:0] Accumulator_1_io_in;
  wire [9:0] Accumulator_1_io_out;
  wire [4:0] Accumulator_1_io_sel;
  wire  Accumulator_1_io_en;
  wire  Accumulator_1_io_reset;
  wire [3:0] _T_657;
  wire [3:0] _T_658;
  wire [3:0] _T_659;
  wire [3:0] _T_660;
  wire [3:0] _T_661;
  wire [3:0] _T_662;
  wire [3:0] _T_663;
  wire [3:0] _T_664;
  reg [5:0] _T_667;
  reg [31:0] _GEN_646;
  reg [5:0] _T_670;
  reg [31:0] _GEN_647;
  reg [5:0] _T_673;
  reg [31:0] _GEN_648;
  reg [5:0] _T_676;
  reg [31:0] _GEN_649;
  reg [5:0] _T_679;
  reg [31:0] _GEN_650;
  reg [5:0] _T_682;
  reg [31:0] _GEN_651;
  reg [5:0] _T_685;
  reg [31:0] _GEN_652;
  reg [5:0] _T_688;
  reg [31:0] _GEN_653;
  reg [5:0] _T_691;
  reg [31:0] _GEN_654;
  reg [5:0] _T_694;
  reg [31:0] _GEN_655;
  reg [5:0] _T_697;
  reg [31:0] _GEN_656;
  reg [5:0] _T_700;
  reg [31:0] _GEN_657;
  reg [5:0] _T_703;
  reg [31:0] _GEN_658;
  reg [5:0] _T_706;
  reg [31:0] _GEN_659;
  reg [5:0] _T_709;
  reg [31:0] _GEN_660;
  reg [5:0] _T_712;
  reg [31:0] _GEN_661;
  wire [5:0] _T_715_0;
  wire [5:0] _T_715_1;
  wire [5:0] _T_715_2;
  wire [5:0] _T_715_3;
  wire [5:0] _T_715_4;
  wire [5:0] _T_715_5;
  wire [5:0] _T_715_6;
  wire [5:0] _T_715_7;
  wire [5:0] _T_715_8;
  wire [5:0] _T_715_9;
  wire [5:0] _T_715_10;
  wire [5:0] _T_715_11;
  wire [5:0] _T_715_12;
  wire [5:0] _T_715_13;
  wire [5:0] _T_715_14;
  wire [5:0] _T_715_15;
  reg [5:0] _T_737;
  reg [31:0] _GEN_662;
  reg [5:0] _T_740;
  reg [31:0] _GEN_663;
  reg [5:0] _T_743;
  reg [31:0] _GEN_664;
  reg [5:0] _T_746;
  reg [31:0] _GEN_665;
  reg [5:0] _T_749;
  reg [31:0] _GEN_666;
  reg [5:0] _T_752;
  reg [31:0] _GEN_667;
  reg [5:0] _T_755;
  reg [31:0] _GEN_668;
  reg [5:0] _T_758;
  reg [31:0] _GEN_669;
  reg [5:0] _T_761;
  reg [31:0] _GEN_670;
  reg [5:0] _T_764;
  reg [31:0] _GEN_671;
  reg [5:0] _T_767;
  reg [31:0] _GEN_672;
  reg [5:0] _T_770;
  reg [31:0] _GEN_673;
  reg [5:0] _T_773;
  reg [31:0] _GEN_674;
  reg [5:0] _T_776;
  reg [31:0] _GEN_675;
  reg [5:0] _T_779;
  reg [31:0] _GEN_676;
  reg [5:0] _T_782;
  reg [31:0] _GEN_677;
  wire [5:0] _T_785_0;
  wire [5:0] _T_785_1;
  wire [5:0] _T_785_2;
  wire [5:0] _T_785_3;
  wire [5:0] _T_785_4;
  wire [5:0] _T_785_5;
  wire [5:0] _T_785_6;
  wire [5:0] _T_785_7;
  wire [5:0] _T_785_8;
  wire [5:0] _T_785_9;
  wire [5:0] _T_785_10;
  wire [5:0] _T_785_11;
  wire [5:0] _T_785_12;
  wire [5:0] _T_785_13;
  wire [5:0] _T_785_14;
  wire [5:0] _T_785_15;
  reg [5:0] _T_807;
  reg [31:0] _GEN_678;
  reg [5:0] _T_810;
  reg [31:0] _GEN_679;
  reg [5:0] _T_813;
  reg [31:0] _GEN_680;
  reg [5:0] _T_816;
  reg [31:0] _GEN_681;
  reg [5:0] _T_819;
  reg [31:0] _GEN_682;
  reg [5:0] _T_822;
  reg [31:0] _GEN_683;
  reg [5:0] _T_825;
  reg [31:0] _GEN_684;
  reg [5:0] _T_828;
  reg [31:0] _GEN_685;
  reg [5:0] _T_831;
  reg [31:0] _GEN_686;
  reg [5:0] _T_834;
  reg [31:0] _GEN_687;
  reg [5:0] _T_837;
  reg [31:0] _GEN_688;
  reg [5:0] _T_840;
  reg [31:0] _GEN_689;
  reg [5:0] _T_843;
  reg [31:0] _GEN_690;
  reg [5:0] _T_846;
  reg [31:0] _GEN_691;
  reg [5:0] _T_849;
  reg [31:0] _GEN_692;
  reg [5:0] _T_852;
  reg [31:0] _GEN_693;
  wire [5:0] _T_855_0;
  wire [5:0] _T_855_1;
  wire [5:0] _T_855_2;
  wire [5:0] _T_855_3;
  wire [5:0] _T_855_4;
  wire [5:0] _T_855_5;
  wire [5:0] _T_855_6;
  wire [5:0] _T_855_7;
  wire [5:0] _T_855_8;
  wire [5:0] _T_855_9;
  wire [5:0] _T_855_10;
  wire [5:0] _T_855_11;
  wire [5:0] _T_855_12;
  wire [5:0] _T_855_13;
  wire [5:0] _T_855_14;
  wire [5:0] _T_855_15;
  reg [5:0] _T_877;
  reg [31:0] _GEN_694;
  reg [5:0] _T_880;
  reg [31:0] _GEN_695;
  reg [5:0] _T_883;
  reg [31:0] _GEN_696;
  reg [5:0] _T_886;
  reg [31:0] _GEN_697;
  reg [5:0] _T_889;
  reg [31:0] _GEN_698;
  reg [5:0] _T_892;
  reg [31:0] _GEN_699;
  reg [5:0] _T_895;
  reg [31:0] _GEN_700;
  reg [5:0] _T_898;
  reg [31:0] _GEN_701;
  reg [5:0] _T_901;
  reg [31:0] _GEN_702;
  reg [5:0] _T_904;
  reg [31:0] _GEN_703;
  reg [5:0] _T_907;
  reg [31:0] _GEN_704;
  reg [5:0] _T_910;
  reg [31:0] _GEN_705;
  reg [5:0] _T_913;
  reg [31:0] _GEN_706;
  reg [5:0] _T_916;
  reg [31:0] _GEN_707;
  reg [5:0] _T_919;
  reg [31:0] _GEN_708;
  reg [5:0] _T_922;
  reg [31:0] _GEN_709;
  wire [5:0] _T_925_0;
  wire [5:0] _T_925_1;
  wire [5:0] _T_925_2;
  wire [5:0] _T_925_3;
  wire [5:0] _T_925_4;
  wire [5:0] _T_925_5;
  wire [5:0] _T_925_6;
  wire [5:0] _T_925_7;
  wire [5:0] _T_925_8;
  wire [5:0] _T_925_9;
  wire [5:0] _T_925_10;
  wire [5:0] _T_925_11;
  wire [5:0] _T_925_12;
  wire [5:0] _T_925_13;
  wire [5:0] _T_925_14;
  wire [5:0] _T_925_15;
  reg [5:0] _T_947;
  reg [31:0] _GEN_710;
  reg [5:0] _T_950;
  reg [31:0] _GEN_711;
  reg [5:0] _T_953;
  reg [31:0] _GEN_712;
  reg [5:0] _T_956;
  reg [31:0] _GEN_713;
  reg [5:0] _T_959;
  reg [31:0] _GEN_714;
  reg [5:0] _T_962;
  reg [31:0] _GEN_715;
  reg [5:0] _T_965;
  reg [31:0] _GEN_716;
  reg [5:0] _T_968;
  reg [31:0] _GEN_717;
  reg [5:0] _T_971;
  reg [31:0] _GEN_718;
  reg [5:0] _T_974;
  reg [31:0] _GEN_719;
  reg [5:0] _T_977;
  reg [31:0] _GEN_720;
  reg [5:0] _T_980;
  reg [31:0] _GEN_721;
  reg [5:0] _T_983;
  reg [31:0] _GEN_722;
  reg [5:0] _T_986;
  reg [31:0] _GEN_723;
  reg [5:0] _T_989;
  reg [31:0] _GEN_724;
  reg [5:0] _T_992;
  reg [31:0] _GEN_725;
  wire [5:0] _T_995_0;
  wire [5:0] _T_995_1;
  wire [5:0] _T_995_2;
  wire [5:0] _T_995_3;
  wire [5:0] _T_995_4;
  wire [5:0] _T_995_5;
  wire [5:0] _T_995_6;
  wire [5:0] _T_995_7;
  wire [5:0] _T_995_8;
  wire [5:0] _T_995_9;
  wire [5:0] _T_995_10;
  wire [5:0] _T_995_11;
  wire [5:0] _T_995_12;
  wire [5:0] _T_995_13;
  wire [5:0] _T_995_14;
  wire [5:0] _T_995_15;
  reg [5:0] _T_1017;
  reg [31:0] _GEN_726;
  reg [5:0] _T_1020;
  reg [31:0] _GEN_727;
  reg [5:0] _T_1023;
  reg [31:0] _GEN_728;
  reg [5:0] _T_1026;
  reg [31:0] _GEN_729;
  reg [5:0] _T_1029;
  reg [31:0] _GEN_730;
  reg [5:0] _T_1032;
  reg [31:0] _GEN_731;
  reg [5:0] _T_1035;
  reg [31:0] _GEN_732;
  reg [5:0] _T_1038;
  reg [31:0] _GEN_733;
  reg [5:0] _T_1041;
  reg [31:0] _GEN_734;
  reg [5:0] _T_1044;
  reg [31:0] _GEN_735;
  reg [5:0] _T_1047;
  reg [31:0] _GEN_736;
  reg [5:0] _T_1050;
  reg [31:0] _GEN_737;
  reg [5:0] _T_1053;
  reg [31:0] _GEN_738;
  reg [5:0] _T_1056;
  reg [31:0] _GEN_739;
  reg [5:0] _T_1059;
  reg [31:0] _GEN_740;
  reg [5:0] _T_1062;
  reg [31:0] _GEN_741;
  wire [5:0] _T_1065_0;
  wire [5:0] _T_1065_1;
  wire [5:0] _T_1065_2;
  wire [5:0] _T_1065_3;
  wire [5:0] _T_1065_4;
  wire [5:0] _T_1065_5;
  wire [5:0] _T_1065_6;
  wire [5:0] _T_1065_7;
  wire [5:0] _T_1065_8;
  wire [5:0] _T_1065_9;
  wire [5:0] _T_1065_10;
  wire [5:0] _T_1065_11;
  wire [5:0] _T_1065_12;
  wire [5:0] _T_1065_13;
  wire [5:0] _T_1065_14;
  wire [5:0] _T_1065_15;
  reg [5:0] _T_1087;
  reg [31:0] _GEN_742;
  reg [5:0] _T_1090;
  reg [31:0] _GEN_743;
  reg [5:0] _T_1093;
  reg [31:0] _GEN_744;
  reg [5:0] _T_1096;
  reg [31:0] _GEN_745;
  reg [5:0] _T_1099;
  reg [31:0] _GEN_746;
  reg [5:0] _T_1102;
  reg [31:0] _GEN_747;
  reg [5:0] _T_1105;
  reg [31:0] _GEN_748;
  reg [5:0] _T_1108;
  reg [31:0] _GEN_749;
  reg [5:0] _T_1111;
  reg [31:0] _GEN_750;
  reg [5:0] _T_1114;
  reg [31:0] _GEN_751;
  reg [5:0] _T_1117;
  reg [31:0] _GEN_752;
  reg [5:0] _T_1120;
  reg [31:0] _GEN_753;
  reg [5:0] _T_1123;
  reg [31:0] _GEN_754;
  reg [5:0] _T_1126;
  reg [31:0] _GEN_755;
  reg [5:0] _T_1129;
  reg [31:0] _GEN_756;
  reg [5:0] _T_1132;
  reg [31:0] _GEN_757;
  wire [5:0] _T_1135_0;
  wire [5:0] _T_1135_1;
  wire [5:0] _T_1135_2;
  wire [5:0] _T_1135_3;
  wire [5:0] _T_1135_4;
  wire [5:0] _T_1135_5;
  wire [5:0] _T_1135_6;
  wire [5:0] _T_1135_7;
  wire [5:0] _T_1135_8;
  wire [5:0] _T_1135_9;
  wire [5:0] _T_1135_10;
  wire [5:0] _T_1135_11;
  wire [5:0] _T_1135_12;
  wire [5:0] _T_1135_13;
  wire [5:0] _T_1135_14;
  wire [5:0] _T_1135_15;
  reg [5:0] _T_1157;
  reg [31:0] _GEN_758;
  reg [5:0] _T_1160;
  reg [31:0] _GEN_759;
  reg [5:0] _T_1163;
  reg [31:0] _GEN_760;
  reg [5:0] _T_1166;
  reg [31:0] _GEN_761;
  reg [5:0] _T_1169;
  reg [31:0] _GEN_762;
  reg [5:0] _T_1172;
  reg [31:0] _GEN_763;
  reg [5:0] _T_1175;
  reg [31:0] _GEN_764;
  reg [5:0] _T_1178;
  reg [31:0] _GEN_765;
  reg [5:0] _T_1181;
  reg [31:0] _GEN_766;
  reg [5:0] _T_1184;
  reg [31:0] _GEN_767;
  reg [5:0] _T_1187;
  reg [31:0] _GEN_768;
  reg [5:0] _T_1190;
  reg [31:0] _GEN_769;
  reg [5:0] _T_1193;
  reg [31:0] _GEN_770;
  reg [5:0] _T_1196;
  reg [31:0] _GEN_771;
  reg [5:0] _T_1199;
  reg [31:0] _GEN_772;
  reg [5:0] _T_1202;
  reg [31:0] _GEN_773;
  wire [5:0] _T_1205_0;
  wire [5:0] _T_1205_1;
  wire [5:0] _T_1205_2;
  wire [5:0] _T_1205_3;
  wire [5:0] _T_1205_4;
  wire [5:0] _T_1205_5;
  wire [5:0] _T_1205_6;
  wire [5:0] _T_1205_7;
  wire [5:0] _T_1205_8;
  wire [5:0] _T_1205_9;
  wire [5:0] _T_1205_10;
  wire [5:0] _T_1205_11;
  wire [5:0] _T_1205_12;
  wire [5:0] _T_1205_13;
  wire [5:0] _T_1205_14;
  wire [5:0] _T_1205_15;
  wire [5:0] _GEN_8;
  wire [5:0] _GEN_152;
  wire [5:0] _GEN_153;
  wire [5:0] _GEN_154;
  wire [5:0] _GEN_155;
  wire [5:0] _GEN_156;
  wire [5:0] _GEN_157;
  wire [5:0] _GEN_158;
  wire [5:0] _GEN_159;
  wire [5:0] _GEN_160;
  wire [5:0] _GEN_161;
  wire [5:0] _GEN_162;
  wire [5:0] _GEN_163;
  wire [5:0] _GEN_164;
  wire [5:0] _GEN_165;
  wire [5:0] _GEN_166;
  wire [5:0] _GEN_9;
  wire [5:0] _GEN_167;
  wire [5:0] _GEN_168;
  wire [5:0] _GEN_169;
  wire [5:0] _GEN_170;
  wire [5:0] _GEN_171;
  wire [5:0] _GEN_172;
  wire [5:0] _GEN_173;
  wire [5:0] _GEN_174;
  wire [5:0] _GEN_175;
  wire [5:0] _GEN_176;
  wire [5:0] _GEN_177;
  wire [5:0] _GEN_178;
  wire [5:0] _GEN_179;
  wire [5:0] _GEN_180;
  wire [5:0] _GEN_181;
  wire [6:0] _T_1225;
  wire [5:0] _T_1226;
  wire [5:0] _T_1227;
  wire [5:0] _GEN_10;
  wire [5:0] _GEN_182;
  wire [5:0] _GEN_183;
  wire [5:0] _GEN_184;
  wire [5:0] _GEN_185;
  wire [5:0] _GEN_186;
  wire [5:0] _GEN_187;
  wire [5:0] _GEN_188;
  wire [5:0] _GEN_189;
  wire [5:0] _GEN_190;
  wire [5:0] _GEN_191;
  wire [5:0] _GEN_192;
  wire [5:0] _GEN_193;
  wire [5:0] _GEN_194;
  wire [5:0] _GEN_195;
  wire [5:0] _GEN_196;
  wire [5:0] _GEN_11;
  wire [5:0] _GEN_197;
  wire [5:0] _GEN_198;
  wire [5:0] _GEN_199;
  wire [5:0] _GEN_200;
  wire [5:0] _GEN_201;
  wire [5:0] _GEN_202;
  wire [5:0] _GEN_203;
  wire [5:0] _GEN_204;
  wire [5:0] _GEN_205;
  wire [5:0] _GEN_206;
  wire [5:0] _GEN_207;
  wire [5:0] _GEN_208;
  wire [5:0] _GEN_209;
  wire [5:0] _GEN_210;
  wire [5:0] _GEN_211;
  wire [6:0] _T_1228;
  wire [5:0] _T_1229;
  wire [5:0] _T_1230;
  wire [5:0] _GEN_12;
  wire [5:0] _GEN_212;
  wire [5:0] _GEN_213;
  wire [5:0] _GEN_214;
  wire [5:0] _GEN_215;
  wire [5:0] _GEN_216;
  wire [5:0] _GEN_217;
  wire [5:0] _GEN_218;
  wire [5:0] _GEN_219;
  wire [5:0] _GEN_220;
  wire [5:0] _GEN_221;
  wire [5:0] _GEN_222;
  wire [5:0] _GEN_223;
  wire [5:0] _GEN_224;
  wire [5:0] _GEN_225;
  wire [5:0] _GEN_226;
  wire [5:0] _GEN_13;
  wire [5:0] _GEN_227;
  wire [5:0] _GEN_228;
  wire [5:0] _GEN_229;
  wire [5:0] _GEN_230;
  wire [5:0] _GEN_231;
  wire [5:0] _GEN_232;
  wire [5:0] _GEN_233;
  wire [5:0] _GEN_234;
  wire [5:0] _GEN_235;
  wire [5:0] _GEN_236;
  wire [5:0] _GEN_237;
  wire [5:0] _GEN_238;
  wire [5:0] _GEN_239;
  wire [5:0] _GEN_240;
  wire [5:0] _GEN_241;
  wire [6:0] _T_1231;
  wire [5:0] _T_1232;
  wire [5:0] _T_1233;
  wire [5:0] _GEN_14;
  wire [5:0] _GEN_242;
  wire [5:0] _GEN_243;
  wire [5:0] _GEN_244;
  wire [5:0] _GEN_245;
  wire [5:0] _GEN_246;
  wire [5:0] _GEN_247;
  wire [5:0] _GEN_248;
  wire [5:0] _GEN_249;
  wire [5:0] _GEN_250;
  wire [5:0] _GEN_251;
  wire [5:0] _GEN_252;
  wire [5:0] _GEN_253;
  wire [5:0] _GEN_254;
  wire [5:0] _GEN_255;
  wire [5:0] _GEN_256;
  wire [5:0] _GEN_15;
  wire [5:0] _GEN_257;
  wire [5:0] _GEN_258;
  wire [5:0] _GEN_259;
  wire [5:0] _GEN_260;
  wire [5:0] _GEN_261;
  wire [5:0] _GEN_262;
  wire [5:0] _GEN_263;
  wire [5:0] _GEN_264;
  wire [5:0] _GEN_265;
  wire [5:0] _GEN_266;
  wire [5:0] _GEN_267;
  wire [5:0] _GEN_268;
  wire [5:0] _GEN_269;
  wire [5:0] _GEN_270;
  wire [5:0] _GEN_271;
  wire [6:0] _T_1234;
  wire [5:0] _T_1235;
  wire [5:0] _T_1236;
  wire [6:0] _T_1237;
  wire [5:0] _T_1238;
  wire [5:0] _T_1239;
  wire [6:0] _T_1240;
  wire [5:0] _T_1241;
  wire [5:0] _T_1242;
  wire [6:0] _T_1243;
  wire [5:0] _T_1244;
  wire [5:0] _T_1245;
  wire [15:0] MulAdd_1_io_a;
  wire [9:0] MulAdd_1_io_b;
  wire [31:0] MulAdd_1_io_m;
  wire [15:0] MulAdd_1_io_c;
  wire [31:0] MulAdd_1_io_r;
  wire [31:0] _T_1246;
  wire [15:0] _T_1247;
  wire [15:0] _T_1248;
  wire [15:0] _T_1249;
  wire [15:0] _T_1250;
  wire  _T_1251;
  wire  signs_1;
  wire  Accumulator_2_clock;
  wire  Accumulator_2_reset;
  wire [9:0] Accumulator_2_io_in;
  wire [9:0] Accumulator_2_io_out;
  wire [4:0] Accumulator_2_io_sel;
  wire  Accumulator_2_io_en;
  wire  Accumulator_2_io_reset;
  wire [3:0] _T_1252;
  wire [3:0] _T_1253;
  wire [3:0] _T_1254;
  wire [3:0] _T_1255;
  wire [3:0] _T_1256;
  wire [3:0] _T_1257;
  wire [3:0] _T_1258;
  wire [3:0] _T_1259;
  reg [5:0] _T_1262;
  reg [31:0] _GEN_774;
  reg [5:0] _T_1265;
  reg [31:0] _GEN_775;
  reg [5:0] _T_1268;
  reg [31:0] _GEN_776;
  reg [5:0] _T_1271;
  reg [31:0] _GEN_777;
  reg [5:0] _T_1274;
  reg [31:0] _GEN_778;
  reg [5:0] _T_1277;
  reg [31:0] _GEN_779;
  reg [5:0] _T_1280;
  reg [31:0] _GEN_780;
  reg [5:0] _T_1283;
  reg [31:0] _GEN_781;
  reg [5:0] _T_1286;
  reg [31:0] _GEN_782;
  reg [5:0] _T_1289;
  reg [31:0] _GEN_783;
  reg [5:0] _T_1292;
  reg [31:0] _GEN_784;
  reg [5:0] _T_1295;
  reg [31:0] _GEN_785;
  reg [5:0] _T_1298;
  reg [31:0] _GEN_786;
  reg [5:0] _T_1301;
  reg [31:0] _GEN_787;
  reg [5:0] _T_1304;
  reg [31:0] _GEN_788;
  reg [5:0] _T_1307;
  reg [31:0] _GEN_789;
  wire [5:0] _T_1310_0;
  wire [5:0] _T_1310_1;
  wire [5:0] _T_1310_2;
  wire [5:0] _T_1310_3;
  wire [5:0] _T_1310_4;
  wire [5:0] _T_1310_5;
  wire [5:0] _T_1310_6;
  wire [5:0] _T_1310_7;
  wire [5:0] _T_1310_8;
  wire [5:0] _T_1310_9;
  wire [5:0] _T_1310_10;
  wire [5:0] _T_1310_11;
  wire [5:0] _T_1310_12;
  wire [5:0] _T_1310_13;
  wire [5:0] _T_1310_14;
  wire [5:0] _T_1310_15;
  reg [5:0] _T_1332;
  reg [31:0] _GEN_790;
  reg [5:0] _T_1335;
  reg [31:0] _GEN_791;
  reg [5:0] _T_1338;
  reg [31:0] _GEN_792;
  reg [5:0] _T_1341;
  reg [31:0] _GEN_793;
  reg [5:0] _T_1344;
  reg [31:0] _GEN_794;
  reg [5:0] _T_1347;
  reg [31:0] _GEN_795;
  reg [5:0] _T_1350;
  reg [31:0] _GEN_796;
  reg [5:0] _T_1353;
  reg [31:0] _GEN_797;
  reg [5:0] _T_1356;
  reg [31:0] _GEN_798;
  reg [5:0] _T_1359;
  reg [31:0] _GEN_799;
  reg [5:0] _T_1362;
  reg [31:0] _GEN_800;
  reg [5:0] _T_1365;
  reg [31:0] _GEN_801;
  reg [5:0] _T_1368;
  reg [31:0] _GEN_802;
  reg [5:0] _T_1371;
  reg [31:0] _GEN_803;
  reg [5:0] _T_1374;
  reg [31:0] _GEN_804;
  reg [5:0] _T_1377;
  reg [31:0] _GEN_805;
  wire [5:0] _T_1380_0;
  wire [5:0] _T_1380_1;
  wire [5:0] _T_1380_2;
  wire [5:0] _T_1380_3;
  wire [5:0] _T_1380_4;
  wire [5:0] _T_1380_5;
  wire [5:0] _T_1380_6;
  wire [5:0] _T_1380_7;
  wire [5:0] _T_1380_8;
  wire [5:0] _T_1380_9;
  wire [5:0] _T_1380_10;
  wire [5:0] _T_1380_11;
  wire [5:0] _T_1380_12;
  wire [5:0] _T_1380_13;
  wire [5:0] _T_1380_14;
  wire [5:0] _T_1380_15;
  reg [5:0] _T_1402;
  reg [31:0] _GEN_806;
  reg [5:0] _T_1405;
  reg [31:0] _GEN_807;
  reg [5:0] _T_1408;
  reg [31:0] _GEN_808;
  reg [5:0] _T_1411;
  reg [31:0] _GEN_809;
  reg [5:0] _T_1414;
  reg [31:0] _GEN_810;
  reg [5:0] _T_1417;
  reg [31:0] _GEN_811;
  reg [5:0] _T_1420;
  reg [31:0] _GEN_812;
  reg [5:0] _T_1423;
  reg [31:0] _GEN_813;
  reg [5:0] _T_1426;
  reg [31:0] _GEN_814;
  reg [5:0] _T_1429;
  reg [31:0] _GEN_815;
  reg [5:0] _T_1432;
  reg [31:0] _GEN_816;
  reg [5:0] _T_1435;
  reg [31:0] _GEN_817;
  reg [5:0] _T_1438;
  reg [31:0] _GEN_818;
  reg [5:0] _T_1441;
  reg [31:0] _GEN_819;
  reg [5:0] _T_1444;
  reg [31:0] _GEN_820;
  reg [5:0] _T_1447;
  reg [31:0] _GEN_821;
  wire [5:0] _T_1450_0;
  wire [5:0] _T_1450_1;
  wire [5:0] _T_1450_2;
  wire [5:0] _T_1450_3;
  wire [5:0] _T_1450_4;
  wire [5:0] _T_1450_5;
  wire [5:0] _T_1450_6;
  wire [5:0] _T_1450_7;
  wire [5:0] _T_1450_8;
  wire [5:0] _T_1450_9;
  wire [5:0] _T_1450_10;
  wire [5:0] _T_1450_11;
  wire [5:0] _T_1450_12;
  wire [5:0] _T_1450_13;
  wire [5:0] _T_1450_14;
  wire [5:0] _T_1450_15;
  reg [5:0] _T_1472;
  reg [31:0] _GEN_822;
  reg [5:0] _T_1475;
  reg [31:0] _GEN_823;
  reg [5:0] _T_1478;
  reg [31:0] _GEN_824;
  reg [5:0] _T_1481;
  reg [31:0] _GEN_825;
  reg [5:0] _T_1484;
  reg [31:0] _GEN_826;
  reg [5:0] _T_1487;
  reg [31:0] _GEN_827;
  reg [5:0] _T_1490;
  reg [31:0] _GEN_828;
  reg [5:0] _T_1493;
  reg [31:0] _GEN_829;
  reg [5:0] _T_1496;
  reg [31:0] _GEN_830;
  reg [5:0] _T_1499;
  reg [31:0] _GEN_831;
  reg [5:0] _T_1502;
  reg [31:0] _GEN_832;
  reg [5:0] _T_1505;
  reg [31:0] _GEN_833;
  reg [5:0] _T_1508;
  reg [31:0] _GEN_834;
  reg [5:0] _T_1511;
  reg [31:0] _GEN_835;
  reg [5:0] _T_1514;
  reg [31:0] _GEN_836;
  reg [5:0] _T_1517;
  reg [31:0] _GEN_837;
  wire [5:0] _T_1520_0;
  wire [5:0] _T_1520_1;
  wire [5:0] _T_1520_2;
  wire [5:0] _T_1520_3;
  wire [5:0] _T_1520_4;
  wire [5:0] _T_1520_5;
  wire [5:0] _T_1520_6;
  wire [5:0] _T_1520_7;
  wire [5:0] _T_1520_8;
  wire [5:0] _T_1520_9;
  wire [5:0] _T_1520_10;
  wire [5:0] _T_1520_11;
  wire [5:0] _T_1520_12;
  wire [5:0] _T_1520_13;
  wire [5:0] _T_1520_14;
  wire [5:0] _T_1520_15;
  reg [5:0] _T_1542;
  reg [31:0] _GEN_838;
  reg [5:0] _T_1545;
  reg [31:0] _GEN_839;
  reg [5:0] _T_1548;
  reg [31:0] _GEN_840;
  reg [5:0] _T_1551;
  reg [31:0] _GEN_841;
  reg [5:0] _T_1554;
  reg [31:0] _GEN_842;
  reg [5:0] _T_1557;
  reg [31:0] _GEN_843;
  reg [5:0] _T_1560;
  reg [31:0] _GEN_844;
  reg [5:0] _T_1563;
  reg [31:0] _GEN_845;
  reg [5:0] _T_1566;
  reg [31:0] _GEN_846;
  reg [5:0] _T_1569;
  reg [31:0] _GEN_847;
  reg [5:0] _T_1572;
  reg [31:0] _GEN_848;
  reg [5:0] _T_1575;
  reg [31:0] _GEN_849;
  reg [5:0] _T_1578;
  reg [31:0] _GEN_850;
  reg [5:0] _T_1581;
  reg [31:0] _GEN_851;
  reg [5:0] _T_1584;
  reg [31:0] _GEN_852;
  reg [5:0] _T_1587;
  reg [31:0] _GEN_853;
  wire [5:0] _T_1590_0;
  wire [5:0] _T_1590_1;
  wire [5:0] _T_1590_2;
  wire [5:0] _T_1590_3;
  wire [5:0] _T_1590_4;
  wire [5:0] _T_1590_5;
  wire [5:0] _T_1590_6;
  wire [5:0] _T_1590_7;
  wire [5:0] _T_1590_8;
  wire [5:0] _T_1590_9;
  wire [5:0] _T_1590_10;
  wire [5:0] _T_1590_11;
  wire [5:0] _T_1590_12;
  wire [5:0] _T_1590_13;
  wire [5:0] _T_1590_14;
  wire [5:0] _T_1590_15;
  reg [5:0] _T_1612;
  reg [31:0] _GEN_854;
  reg [5:0] _T_1615;
  reg [31:0] _GEN_855;
  reg [5:0] _T_1618;
  reg [31:0] _GEN_856;
  reg [5:0] _T_1621;
  reg [31:0] _GEN_857;
  reg [5:0] _T_1624;
  reg [31:0] _GEN_858;
  reg [5:0] _T_1627;
  reg [31:0] _GEN_859;
  reg [5:0] _T_1630;
  reg [31:0] _GEN_860;
  reg [5:0] _T_1633;
  reg [31:0] _GEN_861;
  reg [5:0] _T_1636;
  reg [31:0] _GEN_862;
  reg [5:0] _T_1639;
  reg [31:0] _GEN_863;
  reg [5:0] _T_1642;
  reg [31:0] _GEN_864;
  reg [5:0] _T_1645;
  reg [31:0] _GEN_865;
  reg [5:0] _T_1648;
  reg [31:0] _GEN_866;
  reg [5:0] _T_1651;
  reg [31:0] _GEN_867;
  reg [5:0] _T_1654;
  reg [31:0] _GEN_868;
  reg [5:0] _T_1657;
  reg [31:0] _GEN_869;
  wire [5:0] _T_1660_0;
  wire [5:0] _T_1660_1;
  wire [5:0] _T_1660_2;
  wire [5:0] _T_1660_3;
  wire [5:0] _T_1660_4;
  wire [5:0] _T_1660_5;
  wire [5:0] _T_1660_6;
  wire [5:0] _T_1660_7;
  wire [5:0] _T_1660_8;
  wire [5:0] _T_1660_9;
  wire [5:0] _T_1660_10;
  wire [5:0] _T_1660_11;
  wire [5:0] _T_1660_12;
  wire [5:0] _T_1660_13;
  wire [5:0] _T_1660_14;
  wire [5:0] _T_1660_15;
  reg [5:0] _T_1682;
  reg [31:0] _GEN_870;
  reg [5:0] _T_1685;
  reg [31:0] _GEN_871;
  reg [5:0] _T_1688;
  reg [31:0] _GEN_872;
  reg [5:0] _T_1691;
  reg [31:0] _GEN_873;
  reg [5:0] _T_1694;
  reg [31:0] _GEN_874;
  reg [5:0] _T_1697;
  reg [31:0] _GEN_875;
  reg [5:0] _T_1700;
  reg [31:0] _GEN_876;
  reg [5:0] _T_1703;
  reg [31:0] _GEN_877;
  reg [5:0] _T_1706;
  reg [31:0] _GEN_878;
  reg [5:0] _T_1709;
  reg [31:0] _GEN_879;
  reg [5:0] _T_1712;
  reg [31:0] _GEN_880;
  reg [5:0] _T_1715;
  reg [31:0] _GEN_881;
  reg [5:0] _T_1718;
  reg [31:0] _GEN_882;
  reg [5:0] _T_1721;
  reg [31:0] _GEN_883;
  reg [5:0] _T_1724;
  reg [31:0] _GEN_884;
  reg [5:0] _T_1727;
  reg [31:0] _GEN_885;
  wire [5:0] _T_1730_0;
  wire [5:0] _T_1730_1;
  wire [5:0] _T_1730_2;
  wire [5:0] _T_1730_3;
  wire [5:0] _T_1730_4;
  wire [5:0] _T_1730_5;
  wire [5:0] _T_1730_6;
  wire [5:0] _T_1730_7;
  wire [5:0] _T_1730_8;
  wire [5:0] _T_1730_9;
  wire [5:0] _T_1730_10;
  wire [5:0] _T_1730_11;
  wire [5:0] _T_1730_12;
  wire [5:0] _T_1730_13;
  wire [5:0] _T_1730_14;
  wire [5:0] _T_1730_15;
  reg [5:0] _T_1752;
  reg [31:0] _GEN_886;
  reg [5:0] _T_1755;
  reg [31:0] _GEN_887;
  reg [5:0] _T_1758;
  reg [31:0] _GEN_888;
  reg [5:0] _T_1761;
  reg [31:0] _GEN_889;
  reg [5:0] _T_1764;
  reg [31:0] _GEN_890;
  reg [5:0] _T_1767;
  reg [31:0] _GEN_891;
  reg [5:0] _T_1770;
  reg [31:0] _GEN_892;
  reg [5:0] _T_1773;
  reg [31:0] _GEN_893;
  reg [5:0] _T_1776;
  reg [31:0] _GEN_894;
  reg [5:0] _T_1779;
  reg [31:0] _GEN_895;
  reg [5:0] _T_1782;
  reg [31:0] _GEN_896;
  reg [5:0] _T_1785;
  reg [31:0] _GEN_897;
  reg [5:0] _T_1788;
  reg [31:0] _GEN_898;
  reg [5:0] _T_1791;
  reg [31:0] _GEN_899;
  reg [5:0] _T_1794;
  reg [31:0] _GEN_900;
  reg [5:0] _T_1797;
  reg [31:0] _GEN_901;
  wire [5:0] _T_1800_0;
  wire [5:0] _T_1800_1;
  wire [5:0] _T_1800_2;
  wire [5:0] _T_1800_3;
  wire [5:0] _T_1800_4;
  wire [5:0] _T_1800_5;
  wire [5:0] _T_1800_6;
  wire [5:0] _T_1800_7;
  wire [5:0] _T_1800_8;
  wire [5:0] _T_1800_9;
  wire [5:0] _T_1800_10;
  wire [5:0] _T_1800_11;
  wire [5:0] _T_1800_12;
  wire [5:0] _T_1800_13;
  wire [5:0] _T_1800_14;
  wire [5:0] _T_1800_15;
  wire [5:0] _GEN_16;
  wire [5:0] _GEN_272;
  wire [5:0] _GEN_273;
  wire [5:0] _GEN_274;
  wire [5:0] _GEN_275;
  wire [5:0] _GEN_276;
  wire [5:0] _GEN_277;
  wire [5:0] _GEN_278;
  wire [5:0] _GEN_279;
  wire [5:0] _GEN_280;
  wire [5:0] _GEN_281;
  wire [5:0] _GEN_282;
  wire [5:0] _GEN_283;
  wire [5:0] _GEN_284;
  wire [5:0] _GEN_285;
  wire [5:0] _GEN_286;
  wire [5:0] _GEN_17;
  wire [5:0] _GEN_287;
  wire [5:0] _GEN_288;
  wire [5:0] _GEN_289;
  wire [5:0] _GEN_290;
  wire [5:0] _GEN_291;
  wire [5:0] _GEN_292;
  wire [5:0] _GEN_293;
  wire [5:0] _GEN_294;
  wire [5:0] _GEN_295;
  wire [5:0] _GEN_296;
  wire [5:0] _GEN_297;
  wire [5:0] _GEN_298;
  wire [5:0] _GEN_299;
  wire [5:0] _GEN_300;
  wire [5:0] _GEN_301;
  wire [6:0] _T_1820;
  wire [5:0] _T_1821;
  wire [5:0] _T_1822;
  wire [5:0] _GEN_18;
  wire [5:0] _GEN_302;
  wire [5:0] _GEN_303;
  wire [5:0] _GEN_304;
  wire [5:0] _GEN_305;
  wire [5:0] _GEN_306;
  wire [5:0] _GEN_307;
  wire [5:0] _GEN_308;
  wire [5:0] _GEN_309;
  wire [5:0] _GEN_310;
  wire [5:0] _GEN_311;
  wire [5:0] _GEN_312;
  wire [5:0] _GEN_313;
  wire [5:0] _GEN_314;
  wire [5:0] _GEN_315;
  wire [5:0] _GEN_316;
  wire [5:0] _GEN_19;
  wire [5:0] _GEN_317;
  wire [5:0] _GEN_318;
  wire [5:0] _GEN_319;
  wire [5:0] _GEN_320;
  wire [5:0] _GEN_321;
  wire [5:0] _GEN_322;
  wire [5:0] _GEN_323;
  wire [5:0] _GEN_324;
  wire [5:0] _GEN_325;
  wire [5:0] _GEN_326;
  wire [5:0] _GEN_327;
  wire [5:0] _GEN_328;
  wire [5:0] _GEN_329;
  wire [5:0] _GEN_330;
  wire [5:0] _GEN_331;
  wire [6:0] _T_1823;
  wire [5:0] _T_1824;
  wire [5:0] _T_1825;
  wire [5:0] _GEN_20;
  wire [5:0] _GEN_332;
  wire [5:0] _GEN_333;
  wire [5:0] _GEN_334;
  wire [5:0] _GEN_335;
  wire [5:0] _GEN_336;
  wire [5:0] _GEN_337;
  wire [5:0] _GEN_338;
  wire [5:0] _GEN_339;
  wire [5:0] _GEN_340;
  wire [5:0] _GEN_341;
  wire [5:0] _GEN_342;
  wire [5:0] _GEN_343;
  wire [5:0] _GEN_344;
  wire [5:0] _GEN_345;
  wire [5:0] _GEN_346;
  wire [5:0] _GEN_21;
  wire [5:0] _GEN_347;
  wire [5:0] _GEN_348;
  wire [5:0] _GEN_349;
  wire [5:0] _GEN_350;
  wire [5:0] _GEN_351;
  wire [5:0] _GEN_352;
  wire [5:0] _GEN_353;
  wire [5:0] _GEN_354;
  wire [5:0] _GEN_355;
  wire [5:0] _GEN_356;
  wire [5:0] _GEN_357;
  wire [5:0] _GEN_358;
  wire [5:0] _GEN_359;
  wire [5:0] _GEN_360;
  wire [5:0] _GEN_361;
  wire [6:0] _T_1826;
  wire [5:0] _T_1827;
  wire [5:0] _T_1828;
  wire [5:0] _GEN_22;
  wire [5:0] _GEN_362;
  wire [5:0] _GEN_363;
  wire [5:0] _GEN_364;
  wire [5:0] _GEN_365;
  wire [5:0] _GEN_366;
  wire [5:0] _GEN_367;
  wire [5:0] _GEN_368;
  wire [5:0] _GEN_369;
  wire [5:0] _GEN_370;
  wire [5:0] _GEN_371;
  wire [5:0] _GEN_372;
  wire [5:0] _GEN_373;
  wire [5:0] _GEN_374;
  wire [5:0] _GEN_375;
  wire [5:0] _GEN_376;
  wire [5:0] _GEN_23;
  wire [5:0] _GEN_377;
  wire [5:0] _GEN_378;
  wire [5:0] _GEN_379;
  wire [5:0] _GEN_380;
  wire [5:0] _GEN_381;
  wire [5:0] _GEN_382;
  wire [5:0] _GEN_383;
  wire [5:0] _GEN_384;
  wire [5:0] _GEN_385;
  wire [5:0] _GEN_386;
  wire [5:0] _GEN_387;
  wire [5:0] _GEN_388;
  wire [5:0] _GEN_389;
  wire [5:0] _GEN_390;
  wire [5:0] _GEN_391;
  wire [6:0] _T_1829;
  wire [5:0] _T_1830;
  wire [5:0] _T_1831;
  wire [6:0] _T_1832;
  wire [5:0] _T_1833;
  wire [5:0] _T_1834;
  wire [6:0] _T_1835;
  wire [5:0] _T_1836;
  wire [5:0] _T_1837;
  wire [6:0] _T_1838;
  wire [5:0] _T_1839;
  wire [5:0] _T_1840;
  wire [15:0] MulAdd_2_io_a;
  wire [9:0] MulAdd_2_io_b;
  wire [31:0] MulAdd_2_io_m;
  wire [15:0] MulAdd_2_io_c;
  wire [31:0] MulAdd_2_io_r;
  wire [31:0] _T_1841;
  wire [15:0] _T_1842;
  wire [15:0] _T_1843;
  wire [15:0] _T_1844;
  wire [15:0] _T_1845;
  wire  _T_1846;
  wire  signs_2;
  wire  Accumulator_3_clock;
  wire  Accumulator_3_reset;
  wire [9:0] Accumulator_3_io_in;
  wire [9:0] Accumulator_3_io_out;
  wire [4:0] Accumulator_3_io_sel;
  wire  Accumulator_3_io_en;
  wire  Accumulator_3_io_reset;
  wire [3:0] _T_1847;
  wire [3:0] _T_1848;
  wire [3:0] _T_1849;
  wire [3:0] _T_1850;
  wire [3:0] _T_1851;
  wire [3:0] _T_1852;
  wire [3:0] _T_1853;
  wire [3:0] _T_1854;
  reg [5:0] _T_1857;
  reg [31:0] _GEN_902;
  reg [5:0] _T_1860;
  reg [31:0] _GEN_903;
  reg [5:0] _T_1863;
  reg [31:0] _GEN_904;
  reg [5:0] _T_1866;
  reg [31:0] _GEN_905;
  reg [5:0] _T_1869;
  reg [31:0] _GEN_906;
  reg [5:0] _T_1872;
  reg [31:0] _GEN_907;
  reg [5:0] _T_1875;
  reg [31:0] _GEN_908;
  reg [5:0] _T_1878;
  reg [31:0] _GEN_909;
  reg [5:0] _T_1881;
  reg [31:0] _GEN_910;
  reg [5:0] _T_1884;
  reg [31:0] _GEN_911;
  reg [5:0] _T_1887;
  reg [31:0] _GEN_912;
  reg [5:0] _T_1890;
  reg [31:0] _GEN_913;
  reg [5:0] _T_1893;
  reg [31:0] _GEN_914;
  reg [5:0] _T_1896;
  reg [31:0] _GEN_915;
  reg [5:0] _T_1899;
  reg [31:0] _GEN_916;
  reg [5:0] _T_1902;
  reg [31:0] _GEN_917;
  wire [5:0] _T_1905_0;
  wire [5:0] _T_1905_1;
  wire [5:0] _T_1905_2;
  wire [5:0] _T_1905_3;
  wire [5:0] _T_1905_4;
  wire [5:0] _T_1905_5;
  wire [5:0] _T_1905_6;
  wire [5:0] _T_1905_7;
  wire [5:0] _T_1905_8;
  wire [5:0] _T_1905_9;
  wire [5:0] _T_1905_10;
  wire [5:0] _T_1905_11;
  wire [5:0] _T_1905_12;
  wire [5:0] _T_1905_13;
  wire [5:0] _T_1905_14;
  wire [5:0] _T_1905_15;
  reg [5:0] _T_1927;
  reg [31:0] _GEN_918;
  reg [5:0] _T_1930;
  reg [31:0] _GEN_919;
  reg [5:0] _T_1933;
  reg [31:0] _GEN_920;
  reg [5:0] _T_1936;
  reg [31:0] _GEN_921;
  reg [5:0] _T_1939;
  reg [31:0] _GEN_922;
  reg [5:0] _T_1942;
  reg [31:0] _GEN_923;
  reg [5:0] _T_1945;
  reg [31:0] _GEN_924;
  reg [5:0] _T_1948;
  reg [31:0] _GEN_925;
  reg [5:0] _T_1951;
  reg [31:0] _GEN_926;
  reg [5:0] _T_1954;
  reg [31:0] _GEN_927;
  reg [5:0] _T_1957;
  reg [31:0] _GEN_928;
  reg [5:0] _T_1960;
  reg [31:0] _GEN_929;
  reg [5:0] _T_1963;
  reg [31:0] _GEN_930;
  reg [5:0] _T_1966;
  reg [31:0] _GEN_931;
  reg [5:0] _T_1969;
  reg [31:0] _GEN_932;
  reg [5:0] _T_1972;
  reg [31:0] _GEN_933;
  wire [5:0] _T_1975_0;
  wire [5:0] _T_1975_1;
  wire [5:0] _T_1975_2;
  wire [5:0] _T_1975_3;
  wire [5:0] _T_1975_4;
  wire [5:0] _T_1975_5;
  wire [5:0] _T_1975_6;
  wire [5:0] _T_1975_7;
  wire [5:0] _T_1975_8;
  wire [5:0] _T_1975_9;
  wire [5:0] _T_1975_10;
  wire [5:0] _T_1975_11;
  wire [5:0] _T_1975_12;
  wire [5:0] _T_1975_13;
  wire [5:0] _T_1975_14;
  wire [5:0] _T_1975_15;
  reg [5:0] _T_1997;
  reg [31:0] _GEN_934;
  reg [5:0] _T_2000;
  reg [31:0] _GEN_935;
  reg [5:0] _T_2003;
  reg [31:0] _GEN_936;
  reg [5:0] _T_2006;
  reg [31:0] _GEN_937;
  reg [5:0] _T_2009;
  reg [31:0] _GEN_938;
  reg [5:0] _T_2012;
  reg [31:0] _GEN_939;
  reg [5:0] _T_2015;
  reg [31:0] _GEN_940;
  reg [5:0] _T_2018;
  reg [31:0] _GEN_941;
  reg [5:0] _T_2021;
  reg [31:0] _GEN_942;
  reg [5:0] _T_2024;
  reg [31:0] _GEN_943;
  reg [5:0] _T_2027;
  reg [31:0] _GEN_944;
  reg [5:0] _T_2030;
  reg [31:0] _GEN_945;
  reg [5:0] _T_2033;
  reg [31:0] _GEN_946;
  reg [5:0] _T_2036;
  reg [31:0] _GEN_947;
  reg [5:0] _T_2039;
  reg [31:0] _GEN_948;
  reg [5:0] _T_2042;
  reg [31:0] _GEN_949;
  wire [5:0] _T_2045_0;
  wire [5:0] _T_2045_1;
  wire [5:0] _T_2045_2;
  wire [5:0] _T_2045_3;
  wire [5:0] _T_2045_4;
  wire [5:0] _T_2045_5;
  wire [5:0] _T_2045_6;
  wire [5:0] _T_2045_7;
  wire [5:0] _T_2045_8;
  wire [5:0] _T_2045_9;
  wire [5:0] _T_2045_10;
  wire [5:0] _T_2045_11;
  wire [5:0] _T_2045_12;
  wire [5:0] _T_2045_13;
  wire [5:0] _T_2045_14;
  wire [5:0] _T_2045_15;
  reg [5:0] _T_2067;
  reg [31:0] _GEN_950;
  reg [5:0] _T_2070;
  reg [31:0] _GEN_951;
  reg [5:0] _T_2073;
  reg [31:0] _GEN_952;
  reg [5:0] _T_2076;
  reg [31:0] _GEN_953;
  reg [5:0] _T_2079;
  reg [31:0] _GEN_954;
  reg [5:0] _T_2082;
  reg [31:0] _GEN_955;
  reg [5:0] _T_2085;
  reg [31:0] _GEN_956;
  reg [5:0] _T_2088;
  reg [31:0] _GEN_957;
  reg [5:0] _T_2091;
  reg [31:0] _GEN_958;
  reg [5:0] _T_2094;
  reg [31:0] _GEN_959;
  reg [5:0] _T_2097;
  reg [31:0] _GEN_960;
  reg [5:0] _T_2100;
  reg [31:0] _GEN_961;
  reg [5:0] _T_2103;
  reg [31:0] _GEN_962;
  reg [5:0] _T_2106;
  reg [31:0] _GEN_963;
  reg [5:0] _T_2109;
  reg [31:0] _GEN_964;
  reg [5:0] _T_2112;
  reg [31:0] _GEN_965;
  wire [5:0] _T_2115_0;
  wire [5:0] _T_2115_1;
  wire [5:0] _T_2115_2;
  wire [5:0] _T_2115_3;
  wire [5:0] _T_2115_4;
  wire [5:0] _T_2115_5;
  wire [5:0] _T_2115_6;
  wire [5:0] _T_2115_7;
  wire [5:0] _T_2115_8;
  wire [5:0] _T_2115_9;
  wire [5:0] _T_2115_10;
  wire [5:0] _T_2115_11;
  wire [5:0] _T_2115_12;
  wire [5:0] _T_2115_13;
  wire [5:0] _T_2115_14;
  wire [5:0] _T_2115_15;
  reg [5:0] _T_2137;
  reg [31:0] _GEN_966;
  reg [5:0] _T_2140;
  reg [31:0] _GEN_967;
  reg [5:0] _T_2143;
  reg [31:0] _GEN_968;
  reg [5:0] _T_2146;
  reg [31:0] _GEN_969;
  reg [5:0] _T_2149;
  reg [31:0] _GEN_970;
  reg [5:0] _T_2152;
  reg [31:0] _GEN_971;
  reg [5:0] _T_2155;
  reg [31:0] _GEN_972;
  reg [5:0] _T_2158;
  reg [31:0] _GEN_973;
  reg [5:0] _T_2161;
  reg [31:0] _GEN_974;
  reg [5:0] _T_2164;
  reg [31:0] _GEN_975;
  reg [5:0] _T_2167;
  reg [31:0] _GEN_976;
  reg [5:0] _T_2170;
  reg [31:0] _GEN_977;
  reg [5:0] _T_2173;
  reg [31:0] _GEN_978;
  reg [5:0] _T_2176;
  reg [31:0] _GEN_979;
  reg [5:0] _T_2179;
  reg [31:0] _GEN_980;
  reg [5:0] _T_2182;
  reg [31:0] _GEN_981;
  wire [5:0] _T_2185_0;
  wire [5:0] _T_2185_1;
  wire [5:0] _T_2185_2;
  wire [5:0] _T_2185_3;
  wire [5:0] _T_2185_4;
  wire [5:0] _T_2185_5;
  wire [5:0] _T_2185_6;
  wire [5:0] _T_2185_7;
  wire [5:0] _T_2185_8;
  wire [5:0] _T_2185_9;
  wire [5:0] _T_2185_10;
  wire [5:0] _T_2185_11;
  wire [5:0] _T_2185_12;
  wire [5:0] _T_2185_13;
  wire [5:0] _T_2185_14;
  wire [5:0] _T_2185_15;
  reg [5:0] _T_2207;
  reg [31:0] _GEN_982;
  reg [5:0] _T_2210;
  reg [31:0] _GEN_983;
  reg [5:0] _T_2213;
  reg [31:0] _GEN_984;
  reg [5:0] _T_2216;
  reg [31:0] _GEN_985;
  reg [5:0] _T_2219;
  reg [31:0] _GEN_986;
  reg [5:0] _T_2222;
  reg [31:0] _GEN_987;
  reg [5:0] _T_2225;
  reg [31:0] _GEN_988;
  reg [5:0] _T_2228;
  reg [31:0] _GEN_989;
  reg [5:0] _T_2231;
  reg [31:0] _GEN_990;
  reg [5:0] _T_2234;
  reg [31:0] _GEN_991;
  reg [5:0] _T_2237;
  reg [31:0] _GEN_992;
  reg [5:0] _T_2240;
  reg [31:0] _GEN_993;
  reg [5:0] _T_2243;
  reg [31:0] _GEN_994;
  reg [5:0] _T_2246;
  reg [31:0] _GEN_995;
  reg [5:0] _T_2249;
  reg [31:0] _GEN_996;
  reg [5:0] _T_2252;
  reg [31:0] _GEN_997;
  wire [5:0] _T_2255_0;
  wire [5:0] _T_2255_1;
  wire [5:0] _T_2255_2;
  wire [5:0] _T_2255_3;
  wire [5:0] _T_2255_4;
  wire [5:0] _T_2255_5;
  wire [5:0] _T_2255_6;
  wire [5:0] _T_2255_7;
  wire [5:0] _T_2255_8;
  wire [5:0] _T_2255_9;
  wire [5:0] _T_2255_10;
  wire [5:0] _T_2255_11;
  wire [5:0] _T_2255_12;
  wire [5:0] _T_2255_13;
  wire [5:0] _T_2255_14;
  wire [5:0] _T_2255_15;
  reg [5:0] _T_2277;
  reg [31:0] _GEN_998;
  reg [5:0] _T_2280;
  reg [31:0] _GEN_999;
  reg [5:0] _T_2283;
  reg [31:0] _GEN_1000;
  reg [5:0] _T_2286;
  reg [31:0] _GEN_1001;
  reg [5:0] _T_2289;
  reg [31:0] _GEN_1002;
  reg [5:0] _T_2292;
  reg [31:0] _GEN_1003;
  reg [5:0] _T_2295;
  reg [31:0] _GEN_1004;
  reg [5:0] _T_2298;
  reg [31:0] _GEN_1005;
  reg [5:0] _T_2301;
  reg [31:0] _GEN_1006;
  reg [5:0] _T_2304;
  reg [31:0] _GEN_1007;
  reg [5:0] _T_2307;
  reg [31:0] _GEN_1008;
  reg [5:0] _T_2310;
  reg [31:0] _GEN_1009;
  reg [5:0] _T_2313;
  reg [31:0] _GEN_1010;
  reg [5:0] _T_2316;
  reg [31:0] _GEN_1011;
  reg [5:0] _T_2319;
  reg [31:0] _GEN_1012;
  reg [5:0] _T_2322;
  reg [31:0] _GEN_1013;
  wire [5:0] _T_2325_0;
  wire [5:0] _T_2325_1;
  wire [5:0] _T_2325_2;
  wire [5:0] _T_2325_3;
  wire [5:0] _T_2325_4;
  wire [5:0] _T_2325_5;
  wire [5:0] _T_2325_6;
  wire [5:0] _T_2325_7;
  wire [5:0] _T_2325_8;
  wire [5:0] _T_2325_9;
  wire [5:0] _T_2325_10;
  wire [5:0] _T_2325_11;
  wire [5:0] _T_2325_12;
  wire [5:0] _T_2325_13;
  wire [5:0] _T_2325_14;
  wire [5:0] _T_2325_15;
  reg [5:0] _T_2347;
  reg [31:0] _GEN_1014;
  reg [5:0] _T_2350;
  reg [31:0] _GEN_1015;
  reg [5:0] _T_2353;
  reg [31:0] _GEN_1016;
  reg [5:0] _T_2356;
  reg [31:0] _GEN_1017;
  reg [5:0] _T_2359;
  reg [31:0] _GEN_1018;
  reg [5:0] _T_2362;
  reg [31:0] _GEN_1019;
  reg [5:0] _T_2365;
  reg [31:0] _GEN_1020;
  reg [5:0] _T_2368;
  reg [31:0] _GEN_1021;
  reg [5:0] _T_2371;
  reg [31:0] _GEN_1022;
  reg [5:0] _T_2374;
  reg [31:0] _GEN_1023;
  reg [5:0] _T_2377;
  reg [31:0] _GEN_1024;
  reg [5:0] _T_2380;
  reg [31:0] _GEN_1025;
  reg [5:0] _T_2383;
  reg [31:0] _GEN_1026;
  reg [5:0] _T_2386;
  reg [31:0] _GEN_1027;
  reg [5:0] _T_2389;
  reg [31:0] _GEN_1028;
  reg [5:0] _T_2392;
  reg [31:0] _GEN_1029;
  wire [5:0] _T_2395_0;
  wire [5:0] _T_2395_1;
  wire [5:0] _T_2395_2;
  wire [5:0] _T_2395_3;
  wire [5:0] _T_2395_4;
  wire [5:0] _T_2395_5;
  wire [5:0] _T_2395_6;
  wire [5:0] _T_2395_7;
  wire [5:0] _T_2395_8;
  wire [5:0] _T_2395_9;
  wire [5:0] _T_2395_10;
  wire [5:0] _T_2395_11;
  wire [5:0] _T_2395_12;
  wire [5:0] _T_2395_13;
  wire [5:0] _T_2395_14;
  wire [5:0] _T_2395_15;
  wire [5:0] _GEN_24;
  wire [5:0] _GEN_392;
  wire [5:0] _GEN_393;
  wire [5:0] _GEN_394;
  wire [5:0] _GEN_395;
  wire [5:0] _GEN_396;
  wire [5:0] _GEN_397;
  wire [5:0] _GEN_398;
  wire [5:0] _GEN_399;
  wire [5:0] _GEN_400;
  wire [5:0] _GEN_401;
  wire [5:0] _GEN_402;
  wire [5:0] _GEN_403;
  wire [5:0] _GEN_404;
  wire [5:0] _GEN_405;
  wire [5:0] _GEN_406;
  wire [5:0] _GEN_25;
  wire [5:0] _GEN_407;
  wire [5:0] _GEN_408;
  wire [5:0] _GEN_409;
  wire [5:0] _GEN_410;
  wire [5:0] _GEN_411;
  wire [5:0] _GEN_412;
  wire [5:0] _GEN_413;
  wire [5:0] _GEN_414;
  wire [5:0] _GEN_415;
  wire [5:0] _GEN_416;
  wire [5:0] _GEN_417;
  wire [5:0] _GEN_418;
  wire [5:0] _GEN_419;
  wire [5:0] _GEN_420;
  wire [5:0] _GEN_421;
  wire [6:0] _T_2415;
  wire [5:0] _T_2416;
  wire [5:0] _T_2417;
  wire [5:0] _GEN_26;
  wire [5:0] _GEN_422;
  wire [5:0] _GEN_423;
  wire [5:0] _GEN_424;
  wire [5:0] _GEN_425;
  wire [5:0] _GEN_426;
  wire [5:0] _GEN_427;
  wire [5:0] _GEN_428;
  wire [5:0] _GEN_429;
  wire [5:0] _GEN_430;
  wire [5:0] _GEN_431;
  wire [5:0] _GEN_432;
  wire [5:0] _GEN_433;
  wire [5:0] _GEN_434;
  wire [5:0] _GEN_435;
  wire [5:0] _GEN_436;
  wire [5:0] _GEN_27;
  wire [5:0] _GEN_437;
  wire [5:0] _GEN_438;
  wire [5:0] _GEN_439;
  wire [5:0] _GEN_440;
  wire [5:0] _GEN_441;
  wire [5:0] _GEN_442;
  wire [5:0] _GEN_443;
  wire [5:0] _GEN_444;
  wire [5:0] _GEN_445;
  wire [5:0] _GEN_446;
  wire [5:0] _GEN_447;
  wire [5:0] _GEN_448;
  wire [5:0] _GEN_449;
  wire [5:0] _GEN_450;
  wire [5:0] _GEN_451;
  wire [6:0] _T_2418;
  wire [5:0] _T_2419;
  wire [5:0] _T_2420;
  wire [5:0] _GEN_28;
  wire [5:0] _GEN_452;
  wire [5:0] _GEN_453;
  wire [5:0] _GEN_454;
  wire [5:0] _GEN_455;
  wire [5:0] _GEN_456;
  wire [5:0] _GEN_457;
  wire [5:0] _GEN_458;
  wire [5:0] _GEN_459;
  wire [5:0] _GEN_460;
  wire [5:0] _GEN_461;
  wire [5:0] _GEN_462;
  wire [5:0] _GEN_463;
  wire [5:0] _GEN_464;
  wire [5:0] _GEN_465;
  wire [5:0] _GEN_466;
  wire [5:0] _GEN_29;
  wire [5:0] _GEN_467;
  wire [5:0] _GEN_468;
  wire [5:0] _GEN_469;
  wire [5:0] _GEN_470;
  wire [5:0] _GEN_471;
  wire [5:0] _GEN_472;
  wire [5:0] _GEN_473;
  wire [5:0] _GEN_474;
  wire [5:0] _GEN_475;
  wire [5:0] _GEN_476;
  wire [5:0] _GEN_477;
  wire [5:0] _GEN_478;
  wire [5:0] _GEN_479;
  wire [5:0] _GEN_480;
  wire [5:0] _GEN_481;
  wire [6:0] _T_2421;
  wire [5:0] _T_2422;
  wire [5:0] _T_2423;
  wire [5:0] _GEN_30;
  wire [5:0] _GEN_482;
  wire [5:0] _GEN_483;
  wire [5:0] _GEN_484;
  wire [5:0] _GEN_485;
  wire [5:0] _GEN_486;
  wire [5:0] _GEN_487;
  wire [5:0] _GEN_488;
  wire [5:0] _GEN_489;
  wire [5:0] _GEN_490;
  wire [5:0] _GEN_491;
  wire [5:0] _GEN_492;
  wire [5:0] _GEN_493;
  wire [5:0] _GEN_494;
  wire [5:0] _GEN_495;
  wire [5:0] _GEN_496;
  wire [5:0] _GEN_31;
  wire [5:0] _GEN_497;
  wire [5:0] _GEN_498;
  wire [5:0] _GEN_499;
  wire [5:0] _GEN_500;
  wire [5:0] _GEN_501;
  wire [5:0] _GEN_502;
  wire [5:0] _GEN_503;
  wire [5:0] _GEN_504;
  wire [5:0] _GEN_505;
  wire [5:0] _GEN_506;
  wire [5:0] _GEN_507;
  wire [5:0] _GEN_508;
  wire [5:0] _GEN_509;
  wire [5:0] _GEN_510;
  wire [5:0] _GEN_511;
  wire [6:0] _T_2424;
  wire [5:0] _T_2425;
  wire [5:0] _T_2426;
  wire [6:0] _T_2427;
  wire [5:0] _T_2428;
  wire [5:0] _T_2429;
  wire [6:0] _T_2430;
  wire [5:0] _T_2431;
  wire [5:0] _T_2432;
  wire [6:0] _T_2433;
  wire [5:0] _T_2434;
  wire [5:0] _T_2435;
  wire [15:0] MulAdd_3_io_a;
  wire [9:0] MulAdd_3_io_b;
  wire [31:0] MulAdd_3_io_m;
  wire [15:0] MulAdd_3_io_c;
  wire [31:0] MulAdd_3_io_r;
  wire [31:0] _T_2436;
  wire [15:0] _T_2437;
  wire [15:0] _T_2438;
  wire [15:0] _T_2439;
  wire [15:0] _T_2440;
  wire  _T_2441;
  wire  signs_3;
  wire [1:0] _T_2442;
  wire [1:0] _T_2443;
  wire [3:0] _T_2444;
  reg [31:0] _GEN_512;
  reg [31:0] _GEN_1030;
  reg [31:0] _GEN_513;
  reg [31:0] _GEN_1031;
  reg [15:0] _GEN_514;
  reg [31:0] _GEN_1032;
  reg [15:0] _GEN_515;
  reg [31:0] _GEN_1033;
  reg [31:0] _GEN_516;
  reg [31:0] _GEN_1034;
  reg [15:0] _GEN_517;
  reg [31:0] _GEN_1035;
  AggregateMem mem (
    .clock(mem_clock),
    .io_addr(mem_io_addr),
    .io_waddr(mem_io_waddr),
    .io_in(mem_io_in),
    .io_out(mem_io_out),
    .io_wen(mem_io_wen),
    .io_ren(mem_io_ren)
  );
  BinaryBuffer binaryBuffer (
    .clock(binaryBuffer_clock),
    .io_reset(binaryBuffer_io_reset),
    .io_in(binaryBuffer_io_in),
    .io_fastin(binaryBuffer_io_fastin),
    .io_push(binaryBuffer_io_push),
    .io_fastpush(binaryBuffer_io_fastpush),
    .io_out(binaryBuffer_io_out),
    .io_pop(binaryBuffer_io_pop)
  );
  XNOR xnor$ (
    .io_in1(xnor$_io_in1),
    .io_in2_0(xnor$_io_in2_0),
    .io_in2_1(xnor$_io_in2_1),
    .io_in2_2(xnor$_io_in2_2),
    .io_in2_3(xnor$_io_in2_3),
    .io_out_0(xnor$_io_out_0),
    .io_out_1(xnor$_io_out_1),
    .io_out_2(xnor$_io_out_2),
    .io_out_3(xnor$_io_out_3)
  );
  MeanBuffer meanBuffer (
    .clock(meanBuffer_clock),
    .io_in_0(meanBuffer_io_in_0),
    .io_in_1(meanBuffer_io_in_1),
    .io_in_2(meanBuffer_io_in_2),
    .io_in_3(meanBuffer_io_in_3),
    .io_cntInverse65536(meanBuffer_io_cntInverse65536),
    .io_reset(meanBuffer_io_reset),
    .io_out(meanBuffer_io_out)
  );
  DelayedOutput mean (
    .clock(mean_clock),
    .reset(mean_reset),
    .io_reset(mean_io_reset),
    .io_input(mean_io_input),
    .io_update(mean_io_update),
    .io_output(mean_io_output)
  );
  MaxBuffer maxModule (
    .clock(maxModule_clock),
    .io_reset(maxModule_io_reset),
    .io_en(maxModule_io_en),
    .io_in_0(maxModule_io_in_0),
    .io_in_1(maxModule_io_in_1),
    .io_in_2(maxModule_io_in_2),
    .io_in_3(maxModule_io_in_3),
    .io_offset(maxModule_io_offset),
    .io_out(maxModule_io_out),
    .io_maxLen(maxModule_io_maxLen)
  );
  Accumulator Accumulator (
    .clock(Accumulator_clock),
    .reset(Accumulator_reset),
    .io_in(Accumulator_io_in),
    .io_out(Accumulator_io_out),
    .io_sel(Accumulator_io_sel),
    .io_en(Accumulator_io_en),
    .io_reset(Accumulator_io_reset)
  );
  MulAdd MulAdd (
    .io_a(MulAdd_io_a),
    .io_b(MulAdd_io_b),
    .io_m(MulAdd_io_m),
    .io_c(MulAdd_io_c),
    .io_r(MulAdd_io_r)
  );
  Accumulator Accumulator_1 (
    .clock(Accumulator_1_clock),
    .reset(Accumulator_1_reset),
    .io_in(Accumulator_1_io_in),
    .io_out(Accumulator_1_io_out),
    .io_sel(Accumulator_1_io_sel),
    .io_en(Accumulator_1_io_en),
    .io_reset(Accumulator_1_io_reset)
  );
  MulAdd MulAdd_1 (
    .io_a(MulAdd_1_io_a),
    .io_b(MulAdd_1_io_b),
    .io_m(MulAdd_1_io_m),
    .io_c(MulAdd_1_io_c),
    .io_r(MulAdd_1_io_r)
  );
  Accumulator Accumulator_2 (
    .clock(Accumulator_2_clock),
    .reset(Accumulator_2_reset),
    .io_in(Accumulator_2_io_in),
    .io_out(Accumulator_2_io_out),
    .io_sel(Accumulator_2_io_sel),
    .io_en(Accumulator_2_io_en),
    .io_reset(Accumulator_2_io_reset)
  );
  MulAdd MulAdd_2 (
    .io_a(MulAdd_2_io_a),
    .io_b(MulAdd_2_io_b),
    .io_m(MulAdd_2_io_m),
    .io_c(MulAdd_2_io_c),
    .io_r(MulAdd_2_io_r)
  );
  Accumulator Accumulator_3 (
    .clock(Accumulator_3_clock),
    .reset(Accumulator_3_reset),
    .io_in(Accumulator_3_io_in),
    .io_out(Accumulator_3_io_out),
    .io_sel(Accumulator_3_io_sel),
    .io_en(Accumulator_3_io_en),
    .io_reset(Accumulator_3_io_reset)
  );
  MulAdd MulAdd_3 (
    .io_a(MulAdd_3_io_a),
    .io_b(MulAdd_3_io_b),
    .io_m(MulAdd_3_io_m),
    .io_c(MulAdd_3_io_c),
    .io_r(MulAdd_3_io_r)
  );
  assign io_memOut = mem_io_out;
  assign io_result = maxModule_io_out;
  assign io_mean = mean_io_output;
  assign io_maa = _GEN_514;
  assign io_mab = _GEN_515;
  assign io_mam = _GEN_516;
  assign io_mac = _GEN_517;
  assign mem_clock = clock;
  assign mem_io_addr = io_memAddr;
  assign mem_io_waddr = io_memWAddr;
  assign mem_io_in = io_memIn;
  assign mem_io_wen = io_memWen;
  assign mem_io_ren = 1'h1;
  assign inputWire = _T_2444;
  assign binaryBuffer_clock = clock;
  assign binaryBuffer_io_reset = io_inputBufferReset;
  assign binaryBuffer_io_in = inputWire;
  assign binaryBuffer_io_fastin = io_input;
  assign binaryBuffer_io_push = io_inputBufferPush;
  assign binaryBuffer_io_fastpush = io_inputPush;
  assign binaryBuffer_io_pop = io_inputBufferPop;
  assign xnor$_io_in1 = binaryBuffer_io_out;
  assign xnor$_io_in2_0 = _T_44_0;
  assign xnor$_io_in2_1 = _T_44_1;
  assign xnor$_io_in2_2 = _T_44_2;
  assign xnor$_io_in2_3 = _T_44_3;
  assign _T_33 = mem_io_out;
  assign _T_44_0 = _T_58;
  assign _T_44_1 = _T_59;
  assign _T_44_2 = _T_60;
  assign _T_44_3 = _T_61;
  assign _T_57 = _T_33;
  assign _T_58 = _T_57[31:0];
  assign _T_59 = _T_57[63:32];
  assign _T_60 = _T_57[95:64];
  assign _T_61 = _T_57[127:96];
  assign meanBuffer_clock = clock;
  assign meanBuffer_io_in_0 = MulAdd_io_r;
  assign meanBuffer_io_in_1 = MulAdd_1_io_r;
  assign meanBuffer_io_in_2 = MulAdd_2_io_r;
  assign meanBuffer_io_in_3 = MulAdd_3_io_r;
  assign meanBuffer_io_cntInverse65536 = io_featureNumInverse65536;
  assign meanBuffer_io_reset = io_meanBufferReset;
  assign mean_clock = clock;
  assign mean_reset = reset;
  assign mean_io_reset = io_meanReset;
  assign mean_io_input = meanBuffer_io_out;
  assign mean_io_update = io_meanUpdate;
  assign maxModule_clock = clock;
  assign maxModule_io_reset = io_maxReset;
  assign maxModule_io_en = io_maxEn;
  assign maxModule_io_in_0 = MulAdd_io_r;
  assign maxModule_io_in_1 = MulAdd_1_io_r;
  assign maxModule_io_in_2 = MulAdd_2_io_r;
  assign maxModule_io_in_3 = MulAdd_3_io_r;
  assign maxModule_io_offset = io_maxOffset;
  assign maxModule_io_maxLen = io_actualFeatureNum[3:0];
  assign Accumulator_clock = clock;
  assign Accumulator_reset = reset;
  assign Accumulator_io_in = {{4{_T_650[5]}},_T_650};
  assign Accumulator_io_sel = io_accSel;
  assign Accumulator_io_en = io_accEn;
  assign Accumulator_io_reset = io_accReset;
  assign _T_62 = xnor$_io_out_3[3:0];
  assign _T_63 = xnor$_io_out_3[7:4];
  assign _T_64 = xnor$_io_out_3[11:8];
  assign _T_65 = xnor$_io_out_3[15:12];
  assign _T_66 = xnor$_io_out_3[19:16];
  assign _T_67 = xnor$_io_out_3[23:20];
  assign _T_68 = xnor$_io_out_3[27:24];
  assign _T_69 = xnor$_io_out_3[31:28];
  assign _T_120_0 = _T_72;
  assign _T_120_1 = _T_75;
  assign _T_120_2 = _T_78;
  assign _T_120_3 = _T_81;
  assign _T_120_4 = _T_84;
  assign _T_120_5 = _T_87;
  assign _T_120_6 = _T_90;
  assign _T_120_7 = _T_93;
  assign _T_120_8 = _T_96;
  assign _T_120_9 = _T_99;
  assign _T_120_10 = _T_102;
  assign _T_120_11 = _T_105;
  assign _T_120_12 = _T_108;
  assign _T_120_13 = _T_111;
  assign _T_120_14 = _T_114;
  assign _T_120_15 = _T_117;
  assign _T_190_0 = _T_142;
  assign _T_190_1 = _T_145;
  assign _T_190_2 = _T_148;
  assign _T_190_3 = _T_151;
  assign _T_190_4 = _T_154;
  assign _T_190_5 = _T_157;
  assign _T_190_6 = _T_160;
  assign _T_190_7 = _T_163;
  assign _T_190_8 = _T_166;
  assign _T_190_9 = _T_169;
  assign _T_190_10 = _T_172;
  assign _T_190_11 = _T_175;
  assign _T_190_12 = _T_178;
  assign _T_190_13 = _T_181;
  assign _T_190_14 = _T_184;
  assign _T_190_15 = _T_187;
  assign _T_260_0 = _T_212;
  assign _T_260_1 = _T_215;
  assign _T_260_2 = _T_218;
  assign _T_260_3 = _T_221;
  assign _T_260_4 = _T_224;
  assign _T_260_5 = _T_227;
  assign _T_260_6 = _T_230;
  assign _T_260_7 = _T_233;
  assign _T_260_8 = _T_236;
  assign _T_260_9 = _T_239;
  assign _T_260_10 = _T_242;
  assign _T_260_11 = _T_245;
  assign _T_260_12 = _T_248;
  assign _T_260_13 = _T_251;
  assign _T_260_14 = _T_254;
  assign _T_260_15 = _T_257;
  assign _T_330_0 = _T_282;
  assign _T_330_1 = _T_285;
  assign _T_330_2 = _T_288;
  assign _T_330_3 = _T_291;
  assign _T_330_4 = _T_294;
  assign _T_330_5 = _T_297;
  assign _T_330_6 = _T_300;
  assign _T_330_7 = _T_303;
  assign _T_330_8 = _T_306;
  assign _T_330_9 = _T_309;
  assign _T_330_10 = _T_312;
  assign _T_330_11 = _T_315;
  assign _T_330_12 = _T_318;
  assign _T_330_13 = _T_321;
  assign _T_330_14 = _T_324;
  assign _T_330_15 = _T_327;
  assign _T_400_0 = _T_352;
  assign _T_400_1 = _T_355;
  assign _T_400_2 = _T_358;
  assign _T_400_3 = _T_361;
  assign _T_400_4 = _T_364;
  assign _T_400_5 = _T_367;
  assign _T_400_6 = _T_370;
  assign _T_400_7 = _T_373;
  assign _T_400_8 = _T_376;
  assign _T_400_9 = _T_379;
  assign _T_400_10 = _T_382;
  assign _T_400_11 = _T_385;
  assign _T_400_12 = _T_388;
  assign _T_400_13 = _T_391;
  assign _T_400_14 = _T_394;
  assign _T_400_15 = _T_397;
  assign _T_470_0 = _T_422;
  assign _T_470_1 = _T_425;
  assign _T_470_2 = _T_428;
  assign _T_470_3 = _T_431;
  assign _T_470_4 = _T_434;
  assign _T_470_5 = _T_437;
  assign _T_470_6 = _T_440;
  assign _T_470_7 = _T_443;
  assign _T_470_8 = _T_446;
  assign _T_470_9 = _T_449;
  assign _T_470_10 = _T_452;
  assign _T_470_11 = _T_455;
  assign _T_470_12 = _T_458;
  assign _T_470_13 = _T_461;
  assign _T_470_14 = _T_464;
  assign _T_470_15 = _T_467;
  assign _T_540_0 = _T_492;
  assign _T_540_1 = _T_495;
  assign _T_540_2 = _T_498;
  assign _T_540_3 = _T_501;
  assign _T_540_4 = _T_504;
  assign _T_540_5 = _T_507;
  assign _T_540_6 = _T_510;
  assign _T_540_7 = _T_513;
  assign _T_540_8 = _T_516;
  assign _T_540_9 = _T_519;
  assign _T_540_10 = _T_522;
  assign _T_540_11 = _T_525;
  assign _T_540_12 = _T_528;
  assign _T_540_13 = _T_531;
  assign _T_540_14 = _T_534;
  assign _T_540_15 = _T_537;
  assign _T_610_0 = _T_562;
  assign _T_610_1 = _T_565;
  assign _T_610_2 = _T_568;
  assign _T_610_3 = _T_571;
  assign _T_610_4 = _T_574;
  assign _T_610_5 = _T_577;
  assign _T_610_6 = _T_580;
  assign _T_610_7 = _T_583;
  assign _T_610_8 = _T_586;
  assign _T_610_9 = _T_589;
  assign _T_610_10 = _T_592;
  assign _T_610_11 = _T_595;
  assign _T_610_12 = _T_598;
  assign _T_610_13 = _T_601;
  assign _T_610_14 = _T_604;
  assign _T_610_15 = _T_607;
  assign _GEN_0 = _GEN_46;
  assign _GEN_32 = 4'h1 == _T_62 ? $signed(_T_120_1) : $signed(_T_120_0);
  assign _GEN_33 = 4'h2 == _T_62 ? $signed(_T_120_2) : $signed(_GEN_32);
  assign _GEN_34 = 4'h3 == _T_62 ? $signed(_T_120_3) : $signed(_GEN_33);
  assign _GEN_35 = 4'h4 == _T_62 ? $signed(_T_120_4) : $signed(_GEN_34);
  assign _GEN_36 = 4'h5 == _T_62 ? $signed(_T_120_5) : $signed(_GEN_35);
  assign _GEN_37 = 4'h6 == _T_62 ? $signed(_T_120_6) : $signed(_GEN_36);
  assign _GEN_38 = 4'h7 == _T_62 ? $signed(_T_120_7) : $signed(_GEN_37);
  assign _GEN_39 = 4'h8 == _T_62 ? $signed(_T_120_8) : $signed(_GEN_38);
  assign _GEN_40 = 4'h9 == _T_62 ? $signed(_T_120_9) : $signed(_GEN_39);
  assign _GEN_41 = 4'ha == _T_62 ? $signed(_T_120_10) : $signed(_GEN_40);
  assign _GEN_42 = 4'hb == _T_62 ? $signed(_T_120_11) : $signed(_GEN_41);
  assign _GEN_43 = 4'hc == _T_62 ? $signed(_T_120_12) : $signed(_GEN_42);
  assign _GEN_44 = 4'hd == _T_62 ? $signed(_T_120_13) : $signed(_GEN_43);
  assign _GEN_45 = 4'he == _T_62 ? $signed(_T_120_14) : $signed(_GEN_44);
  assign _GEN_46 = 4'hf == _T_62 ? $signed(_T_120_15) : $signed(_GEN_45);
  assign _GEN_1 = _GEN_61;
  assign _GEN_47 = 4'h1 == _T_63 ? $signed(_T_190_1) : $signed(_T_190_0);
  assign _GEN_48 = 4'h2 == _T_63 ? $signed(_T_190_2) : $signed(_GEN_47);
  assign _GEN_49 = 4'h3 == _T_63 ? $signed(_T_190_3) : $signed(_GEN_48);
  assign _GEN_50 = 4'h4 == _T_63 ? $signed(_T_190_4) : $signed(_GEN_49);
  assign _GEN_51 = 4'h5 == _T_63 ? $signed(_T_190_5) : $signed(_GEN_50);
  assign _GEN_52 = 4'h6 == _T_63 ? $signed(_T_190_6) : $signed(_GEN_51);
  assign _GEN_53 = 4'h7 == _T_63 ? $signed(_T_190_7) : $signed(_GEN_52);
  assign _GEN_54 = 4'h8 == _T_63 ? $signed(_T_190_8) : $signed(_GEN_53);
  assign _GEN_55 = 4'h9 == _T_63 ? $signed(_T_190_9) : $signed(_GEN_54);
  assign _GEN_56 = 4'ha == _T_63 ? $signed(_T_190_10) : $signed(_GEN_55);
  assign _GEN_57 = 4'hb == _T_63 ? $signed(_T_190_11) : $signed(_GEN_56);
  assign _GEN_58 = 4'hc == _T_63 ? $signed(_T_190_12) : $signed(_GEN_57);
  assign _GEN_59 = 4'hd == _T_63 ? $signed(_T_190_13) : $signed(_GEN_58);
  assign _GEN_60 = 4'he == _T_63 ? $signed(_T_190_14) : $signed(_GEN_59);
  assign _GEN_61 = 4'hf == _T_63 ? $signed(_T_190_15) : $signed(_GEN_60);
  assign _T_630 = $signed(_GEN_0) + $signed(_GEN_1);
  assign _T_631 = _T_630[5:0];
  assign _T_632 = $signed(_T_631);
  assign _GEN_2 = _GEN_76;
  assign _GEN_62 = 4'h1 == _T_64 ? $signed(_T_260_1) : $signed(_T_260_0);
  assign _GEN_63 = 4'h2 == _T_64 ? $signed(_T_260_2) : $signed(_GEN_62);
  assign _GEN_64 = 4'h3 == _T_64 ? $signed(_T_260_3) : $signed(_GEN_63);
  assign _GEN_65 = 4'h4 == _T_64 ? $signed(_T_260_4) : $signed(_GEN_64);
  assign _GEN_66 = 4'h5 == _T_64 ? $signed(_T_260_5) : $signed(_GEN_65);
  assign _GEN_67 = 4'h6 == _T_64 ? $signed(_T_260_6) : $signed(_GEN_66);
  assign _GEN_68 = 4'h7 == _T_64 ? $signed(_T_260_7) : $signed(_GEN_67);
  assign _GEN_69 = 4'h8 == _T_64 ? $signed(_T_260_8) : $signed(_GEN_68);
  assign _GEN_70 = 4'h9 == _T_64 ? $signed(_T_260_9) : $signed(_GEN_69);
  assign _GEN_71 = 4'ha == _T_64 ? $signed(_T_260_10) : $signed(_GEN_70);
  assign _GEN_72 = 4'hb == _T_64 ? $signed(_T_260_11) : $signed(_GEN_71);
  assign _GEN_73 = 4'hc == _T_64 ? $signed(_T_260_12) : $signed(_GEN_72);
  assign _GEN_74 = 4'hd == _T_64 ? $signed(_T_260_13) : $signed(_GEN_73);
  assign _GEN_75 = 4'he == _T_64 ? $signed(_T_260_14) : $signed(_GEN_74);
  assign _GEN_76 = 4'hf == _T_64 ? $signed(_T_260_15) : $signed(_GEN_75);
  assign _GEN_3 = _GEN_91;
  assign _GEN_77 = 4'h1 == _T_65 ? $signed(_T_330_1) : $signed(_T_330_0);
  assign _GEN_78 = 4'h2 == _T_65 ? $signed(_T_330_2) : $signed(_GEN_77);
  assign _GEN_79 = 4'h3 == _T_65 ? $signed(_T_330_3) : $signed(_GEN_78);
  assign _GEN_80 = 4'h4 == _T_65 ? $signed(_T_330_4) : $signed(_GEN_79);
  assign _GEN_81 = 4'h5 == _T_65 ? $signed(_T_330_5) : $signed(_GEN_80);
  assign _GEN_82 = 4'h6 == _T_65 ? $signed(_T_330_6) : $signed(_GEN_81);
  assign _GEN_83 = 4'h7 == _T_65 ? $signed(_T_330_7) : $signed(_GEN_82);
  assign _GEN_84 = 4'h8 == _T_65 ? $signed(_T_330_8) : $signed(_GEN_83);
  assign _GEN_85 = 4'h9 == _T_65 ? $signed(_T_330_9) : $signed(_GEN_84);
  assign _GEN_86 = 4'ha == _T_65 ? $signed(_T_330_10) : $signed(_GEN_85);
  assign _GEN_87 = 4'hb == _T_65 ? $signed(_T_330_11) : $signed(_GEN_86);
  assign _GEN_88 = 4'hc == _T_65 ? $signed(_T_330_12) : $signed(_GEN_87);
  assign _GEN_89 = 4'hd == _T_65 ? $signed(_T_330_13) : $signed(_GEN_88);
  assign _GEN_90 = 4'he == _T_65 ? $signed(_T_330_14) : $signed(_GEN_89);
  assign _GEN_91 = 4'hf == _T_65 ? $signed(_T_330_15) : $signed(_GEN_90);
  assign _T_633 = $signed(_GEN_2) + $signed(_GEN_3);
  assign _T_634 = _T_633[5:0];
  assign _T_635 = $signed(_T_634);
  assign _GEN_4 = _GEN_106;
  assign _GEN_92 = 4'h1 == _T_66 ? $signed(_T_400_1) : $signed(_T_400_0);
  assign _GEN_93 = 4'h2 == _T_66 ? $signed(_T_400_2) : $signed(_GEN_92);
  assign _GEN_94 = 4'h3 == _T_66 ? $signed(_T_400_3) : $signed(_GEN_93);
  assign _GEN_95 = 4'h4 == _T_66 ? $signed(_T_400_4) : $signed(_GEN_94);
  assign _GEN_96 = 4'h5 == _T_66 ? $signed(_T_400_5) : $signed(_GEN_95);
  assign _GEN_97 = 4'h6 == _T_66 ? $signed(_T_400_6) : $signed(_GEN_96);
  assign _GEN_98 = 4'h7 == _T_66 ? $signed(_T_400_7) : $signed(_GEN_97);
  assign _GEN_99 = 4'h8 == _T_66 ? $signed(_T_400_8) : $signed(_GEN_98);
  assign _GEN_100 = 4'h9 == _T_66 ? $signed(_T_400_9) : $signed(_GEN_99);
  assign _GEN_101 = 4'ha == _T_66 ? $signed(_T_400_10) : $signed(_GEN_100);
  assign _GEN_102 = 4'hb == _T_66 ? $signed(_T_400_11) : $signed(_GEN_101);
  assign _GEN_103 = 4'hc == _T_66 ? $signed(_T_400_12) : $signed(_GEN_102);
  assign _GEN_104 = 4'hd == _T_66 ? $signed(_T_400_13) : $signed(_GEN_103);
  assign _GEN_105 = 4'he == _T_66 ? $signed(_T_400_14) : $signed(_GEN_104);
  assign _GEN_106 = 4'hf == _T_66 ? $signed(_T_400_15) : $signed(_GEN_105);
  assign _GEN_5 = _GEN_121;
  assign _GEN_107 = 4'h1 == _T_67 ? $signed(_T_470_1) : $signed(_T_470_0);
  assign _GEN_108 = 4'h2 == _T_67 ? $signed(_T_470_2) : $signed(_GEN_107);
  assign _GEN_109 = 4'h3 == _T_67 ? $signed(_T_470_3) : $signed(_GEN_108);
  assign _GEN_110 = 4'h4 == _T_67 ? $signed(_T_470_4) : $signed(_GEN_109);
  assign _GEN_111 = 4'h5 == _T_67 ? $signed(_T_470_5) : $signed(_GEN_110);
  assign _GEN_112 = 4'h6 == _T_67 ? $signed(_T_470_6) : $signed(_GEN_111);
  assign _GEN_113 = 4'h7 == _T_67 ? $signed(_T_470_7) : $signed(_GEN_112);
  assign _GEN_114 = 4'h8 == _T_67 ? $signed(_T_470_8) : $signed(_GEN_113);
  assign _GEN_115 = 4'h9 == _T_67 ? $signed(_T_470_9) : $signed(_GEN_114);
  assign _GEN_116 = 4'ha == _T_67 ? $signed(_T_470_10) : $signed(_GEN_115);
  assign _GEN_117 = 4'hb == _T_67 ? $signed(_T_470_11) : $signed(_GEN_116);
  assign _GEN_118 = 4'hc == _T_67 ? $signed(_T_470_12) : $signed(_GEN_117);
  assign _GEN_119 = 4'hd == _T_67 ? $signed(_T_470_13) : $signed(_GEN_118);
  assign _GEN_120 = 4'he == _T_67 ? $signed(_T_470_14) : $signed(_GEN_119);
  assign _GEN_121 = 4'hf == _T_67 ? $signed(_T_470_15) : $signed(_GEN_120);
  assign _T_636 = $signed(_GEN_4) + $signed(_GEN_5);
  assign _T_637 = _T_636[5:0];
  assign _T_638 = $signed(_T_637);
  assign _GEN_6 = _GEN_136;
  assign _GEN_122 = 4'h1 == _T_68 ? $signed(_T_540_1) : $signed(_T_540_0);
  assign _GEN_123 = 4'h2 == _T_68 ? $signed(_T_540_2) : $signed(_GEN_122);
  assign _GEN_124 = 4'h3 == _T_68 ? $signed(_T_540_3) : $signed(_GEN_123);
  assign _GEN_125 = 4'h4 == _T_68 ? $signed(_T_540_4) : $signed(_GEN_124);
  assign _GEN_126 = 4'h5 == _T_68 ? $signed(_T_540_5) : $signed(_GEN_125);
  assign _GEN_127 = 4'h6 == _T_68 ? $signed(_T_540_6) : $signed(_GEN_126);
  assign _GEN_128 = 4'h7 == _T_68 ? $signed(_T_540_7) : $signed(_GEN_127);
  assign _GEN_129 = 4'h8 == _T_68 ? $signed(_T_540_8) : $signed(_GEN_128);
  assign _GEN_130 = 4'h9 == _T_68 ? $signed(_T_540_9) : $signed(_GEN_129);
  assign _GEN_131 = 4'ha == _T_68 ? $signed(_T_540_10) : $signed(_GEN_130);
  assign _GEN_132 = 4'hb == _T_68 ? $signed(_T_540_11) : $signed(_GEN_131);
  assign _GEN_133 = 4'hc == _T_68 ? $signed(_T_540_12) : $signed(_GEN_132);
  assign _GEN_134 = 4'hd == _T_68 ? $signed(_T_540_13) : $signed(_GEN_133);
  assign _GEN_135 = 4'he == _T_68 ? $signed(_T_540_14) : $signed(_GEN_134);
  assign _GEN_136 = 4'hf == _T_68 ? $signed(_T_540_15) : $signed(_GEN_135);
  assign _GEN_7 = _GEN_151;
  assign _GEN_137 = 4'h1 == _T_69 ? $signed(_T_610_1) : $signed(_T_610_0);
  assign _GEN_138 = 4'h2 == _T_69 ? $signed(_T_610_2) : $signed(_GEN_137);
  assign _GEN_139 = 4'h3 == _T_69 ? $signed(_T_610_3) : $signed(_GEN_138);
  assign _GEN_140 = 4'h4 == _T_69 ? $signed(_T_610_4) : $signed(_GEN_139);
  assign _GEN_141 = 4'h5 == _T_69 ? $signed(_T_610_5) : $signed(_GEN_140);
  assign _GEN_142 = 4'h6 == _T_69 ? $signed(_T_610_6) : $signed(_GEN_141);
  assign _GEN_143 = 4'h7 == _T_69 ? $signed(_T_610_7) : $signed(_GEN_142);
  assign _GEN_144 = 4'h8 == _T_69 ? $signed(_T_610_8) : $signed(_GEN_143);
  assign _GEN_145 = 4'h9 == _T_69 ? $signed(_T_610_9) : $signed(_GEN_144);
  assign _GEN_146 = 4'ha == _T_69 ? $signed(_T_610_10) : $signed(_GEN_145);
  assign _GEN_147 = 4'hb == _T_69 ? $signed(_T_610_11) : $signed(_GEN_146);
  assign _GEN_148 = 4'hc == _T_69 ? $signed(_T_610_12) : $signed(_GEN_147);
  assign _GEN_149 = 4'hd == _T_69 ? $signed(_T_610_13) : $signed(_GEN_148);
  assign _GEN_150 = 4'he == _T_69 ? $signed(_T_610_14) : $signed(_GEN_149);
  assign _GEN_151 = 4'hf == _T_69 ? $signed(_T_610_15) : $signed(_GEN_150);
  assign _T_639 = $signed(_GEN_6) + $signed(_GEN_7);
  assign _T_640 = _T_639[5:0];
  assign _T_641 = $signed(_T_640);
  assign _T_642 = $signed(_T_632) + $signed(_T_635);
  assign _T_643 = _T_642[5:0];
  assign _T_644 = $signed(_T_643);
  assign _T_645 = $signed(_T_638) + $signed(_T_641);
  assign _T_646 = _T_645[5:0];
  assign _T_647 = $signed(_T_646);
  assign _T_648 = $signed(_T_644) + $signed(_T_647);
  assign _T_649 = _T_648[5:0];
  assign _T_650 = $signed(_T_649);
  assign MulAdd_io_a = _T_653;
  assign MulAdd_io_b = Accumulator_io_out;
  assign MulAdd_io_m = mean_io_output;
  assign MulAdd_io_c = _T_655;
  assign _T_651 = mem_io_out[127:96];
  assign _T_652 = _T_651[31:16];
  assign _T_653 = $signed(_T_652);
  assign _T_654 = _T_651[15:0];
  assign _T_655 = $signed(_T_654);
  assign _T_656 = MulAdd_io_r[31];
  assign signs_0 = ~ _T_656;
  assign Accumulator_1_clock = clock;
  assign Accumulator_1_reset = reset;
  assign Accumulator_1_io_in = {{4{_T_1245[5]}},_T_1245};
  assign Accumulator_1_io_sel = io_accSel;
  assign Accumulator_1_io_en = io_accEn;
  assign Accumulator_1_io_reset = io_accReset;
  assign _T_657 = xnor$_io_out_2[3:0];
  assign _T_658 = xnor$_io_out_2[7:4];
  assign _T_659 = xnor$_io_out_2[11:8];
  assign _T_660 = xnor$_io_out_2[15:12];
  assign _T_661 = xnor$_io_out_2[19:16];
  assign _T_662 = xnor$_io_out_2[23:20];
  assign _T_663 = xnor$_io_out_2[27:24];
  assign _T_664 = xnor$_io_out_2[31:28];
  assign _T_715_0 = _T_667;
  assign _T_715_1 = _T_670;
  assign _T_715_2 = _T_673;
  assign _T_715_3 = _T_676;
  assign _T_715_4 = _T_679;
  assign _T_715_5 = _T_682;
  assign _T_715_6 = _T_685;
  assign _T_715_7 = _T_688;
  assign _T_715_8 = _T_691;
  assign _T_715_9 = _T_694;
  assign _T_715_10 = _T_697;
  assign _T_715_11 = _T_700;
  assign _T_715_12 = _T_703;
  assign _T_715_13 = _T_706;
  assign _T_715_14 = _T_709;
  assign _T_715_15 = _T_712;
  assign _T_785_0 = _T_737;
  assign _T_785_1 = _T_740;
  assign _T_785_2 = _T_743;
  assign _T_785_3 = _T_746;
  assign _T_785_4 = _T_749;
  assign _T_785_5 = _T_752;
  assign _T_785_6 = _T_755;
  assign _T_785_7 = _T_758;
  assign _T_785_8 = _T_761;
  assign _T_785_9 = _T_764;
  assign _T_785_10 = _T_767;
  assign _T_785_11 = _T_770;
  assign _T_785_12 = _T_773;
  assign _T_785_13 = _T_776;
  assign _T_785_14 = _T_779;
  assign _T_785_15 = _T_782;
  assign _T_855_0 = _T_807;
  assign _T_855_1 = _T_810;
  assign _T_855_2 = _T_813;
  assign _T_855_3 = _T_816;
  assign _T_855_4 = _T_819;
  assign _T_855_5 = _T_822;
  assign _T_855_6 = _T_825;
  assign _T_855_7 = _T_828;
  assign _T_855_8 = _T_831;
  assign _T_855_9 = _T_834;
  assign _T_855_10 = _T_837;
  assign _T_855_11 = _T_840;
  assign _T_855_12 = _T_843;
  assign _T_855_13 = _T_846;
  assign _T_855_14 = _T_849;
  assign _T_855_15 = _T_852;
  assign _T_925_0 = _T_877;
  assign _T_925_1 = _T_880;
  assign _T_925_2 = _T_883;
  assign _T_925_3 = _T_886;
  assign _T_925_4 = _T_889;
  assign _T_925_5 = _T_892;
  assign _T_925_6 = _T_895;
  assign _T_925_7 = _T_898;
  assign _T_925_8 = _T_901;
  assign _T_925_9 = _T_904;
  assign _T_925_10 = _T_907;
  assign _T_925_11 = _T_910;
  assign _T_925_12 = _T_913;
  assign _T_925_13 = _T_916;
  assign _T_925_14 = _T_919;
  assign _T_925_15 = _T_922;
  assign _T_995_0 = _T_947;
  assign _T_995_1 = _T_950;
  assign _T_995_2 = _T_953;
  assign _T_995_3 = _T_956;
  assign _T_995_4 = _T_959;
  assign _T_995_5 = _T_962;
  assign _T_995_6 = _T_965;
  assign _T_995_7 = _T_968;
  assign _T_995_8 = _T_971;
  assign _T_995_9 = _T_974;
  assign _T_995_10 = _T_977;
  assign _T_995_11 = _T_980;
  assign _T_995_12 = _T_983;
  assign _T_995_13 = _T_986;
  assign _T_995_14 = _T_989;
  assign _T_995_15 = _T_992;
  assign _T_1065_0 = _T_1017;
  assign _T_1065_1 = _T_1020;
  assign _T_1065_2 = _T_1023;
  assign _T_1065_3 = _T_1026;
  assign _T_1065_4 = _T_1029;
  assign _T_1065_5 = _T_1032;
  assign _T_1065_6 = _T_1035;
  assign _T_1065_7 = _T_1038;
  assign _T_1065_8 = _T_1041;
  assign _T_1065_9 = _T_1044;
  assign _T_1065_10 = _T_1047;
  assign _T_1065_11 = _T_1050;
  assign _T_1065_12 = _T_1053;
  assign _T_1065_13 = _T_1056;
  assign _T_1065_14 = _T_1059;
  assign _T_1065_15 = _T_1062;
  assign _T_1135_0 = _T_1087;
  assign _T_1135_1 = _T_1090;
  assign _T_1135_2 = _T_1093;
  assign _T_1135_3 = _T_1096;
  assign _T_1135_4 = _T_1099;
  assign _T_1135_5 = _T_1102;
  assign _T_1135_6 = _T_1105;
  assign _T_1135_7 = _T_1108;
  assign _T_1135_8 = _T_1111;
  assign _T_1135_9 = _T_1114;
  assign _T_1135_10 = _T_1117;
  assign _T_1135_11 = _T_1120;
  assign _T_1135_12 = _T_1123;
  assign _T_1135_13 = _T_1126;
  assign _T_1135_14 = _T_1129;
  assign _T_1135_15 = _T_1132;
  assign _T_1205_0 = _T_1157;
  assign _T_1205_1 = _T_1160;
  assign _T_1205_2 = _T_1163;
  assign _T_1205_3 = _T_1166;
  assign _T_1205_4 = _T_1169;
  assign _T_1205_5 = _T_1172;
  assign _T_1205_6 = _T_1175;
  assign _T_1205_7 = _T_1178;
  assign _T_1205_8 = _T_1181;
  assign _T_1205_9 = _T_1184;
  assign _T_1205_10 = _T_1187;
  assign _T_1205_11 = _T_1190;
  assign _T_1205_12 = _T_1193;
  assign _T_1205_13 = _T_1196;
  assign _T_1205_14 = _T_1199;
  assign _T_1205_15 = _T_1202;
  assign _GEN_8 = _GEN_166;
  assign _GEN_152 = 4'h1 == _T_657 ? $signed(_T_715_1) : $signed(_T_715_0);
  assign _GEN_153 = 4'h2 == _T_657 ? $signed(_T_715_2) : $signed(_GEN_152);
  assign _GEN_154 = 4'h3 == _T_657 ? $signed(_T_715_3) : $signed(_GEN_153);
  assign _GEN_155 = 4'h4 == _T_657 ? $signed(_T_715_4) : $signed(_GEN_154);
  assign _GEN_156 = 4'h5 == _T_657 ? $signed(_T_715_5) : $signed(_GEN_155);
  assign _GEN_157 = 4'h6 == _T_657 ? $signed(_T_715_6) : $signed(_GEN_156);
  assign _GEN_158 = 4'h7 == _T_657 ? $signed(_T_715_7) : $signed(_GEN_157);
  assign _GEN_159 = 4'h8 == _T_657 ? $signed(_T_715_8) : $signed(_GEN_158);
  assign _GEN_160 = 4'h9 == _T_657 ? $signed(_T_715_9) : $signed(_GEN_159);
  assign _GEN_161 = 4'ha == _T_657 ? $signed(_T_715_10) : $signed(_GEN_160);
  assign _GEN_162 = 4'hb == _T_657 ? $signed(_T_715_11) : $signed(_GEN_161);
  assign _GEN_163 = 4'hc == _T_657 ? $signed(_T_715_12) : $signed(_GEN_162);
  assign _GEN_164 = 4'hd == _T_657 ? $signed(_T_715_13) : $signed(_GEN_163);
  assign _GEN_165 = 4'he == _T_657 ? $signed(_T_715_14) : $signed(_GEN_164);
  assign _GEN_166 = 4'hf == _T_657 ? $signed(_T_715_15) : $signed(_GEN_165);
  assign _GEN_9 = _GEN_181;
  assign _GEN_167 = 4'h1 == _T_658 ? $signed(_T_785_1) : $signed(_T_785_0);
  assign _GEN_168 = 4'h2 == _T_658 ? $signed(_T_785_2) : $signed(_GEN_167);
  assign _GEN_169 = 4'h3 == _T_658 ? $signed(_T_785_3) : $signed(_GEN_168);
  assign _GEN_170 = 4'h4 == _T_658 ? $signed(_T_785_4) : $signed(_GEN_169);
  assign _GEN_171 = 4'h5 == _T_658 ? $signed(_T_785_5) : $signed(_GEN_170);
  assign _GEN_172 = 4'h6 == _T_658 ? $signed(_T_785_6) : $signed(_GEN_171);
  assign _GEN_173 = 4'h7 == _T_658 ? $signed(_T_785_7) : $signed(_GEN_172);
  assign _GEN_174 = 4'h8 == _T_658 ? $signed(_T_785_8) : $signed(_GEN_173);
  assign _GEN_175 = 4'h9 == _T_658 ? $signed(_T_785_9) : $signed(_GEN_174);
  assign _GEN_176 = 4'ha == _T_658 ? $signed(_T_785_10) : $signed(_GEN_175);
  assign _GEN_177 = 4'hb == _T_658 ? $signed(_T_785_11) : $signed(_GEN_176);
  assign _GEN_178 = 4'hc == _T_658 ? $signed(_T_785_12) : $signed(_GEN_177);
  assign _GEN_179 = 4'hd == _T_658 ? $signed(_T_785_13) : $signed(_GEN_178);
  assign _GEN_180 = 4'he == _T_658 ? $signed(_T_785_14) : $signed(_GEN_179);
  assign _GEN_181 = 4'hf == _T_658 ? $signed(_T_785_15) : $signed(_GEN_180);
  assign _T_1225 = $signed(_GEN_8) + $signed(_GEN_9);
  assign _T_1226 = _T_1225[5:0];
  assign _T_1227 = $signed(_T_1226);
  assign _GEN_10 = _GEN_196;
  assign _GEN_182 = 4'h1 == _T_659 ? $signed(_T_855_1) : $signed(_T_855_0);
  assign _GEN_183 = 4'h2 == _T_659 ? $signed(_T_855_2) : $signed(_GEN_182);
  assign _GEN_184 = 4'h3 == _T_659 ? $signed(_T_855_3) : $signed(_GEN_183);
  assign _GEN_185 = 4'h4 == _T_659 ? $signed(_T_855_4) : $signed(_GEN_184);
  assign _GEN_186 = 4'h5 == _T_659 ? $signed(_T_855_5) : $signed(_GEN_185);
  assign _GEN_187 = 4'h6 == _T_659 ? $signed(_T_855_6) : $signed(_GEN_186);
  assign _GEN_188 = 4'h7 == _T_659 ? $signed(_T_855_7) : $signed(_GEN_187);
  assign _GEN_189 = 4'h8 == _T_659 ? $signed(_T_855_8) : $signed(_GEN_188);
  assign _GEN_190 = 4'h9 == _T_659 ? $signed(_T_855_9) : $signed(_GEN_189);
  assign _GEN_191 = 4'ha == _T_659 ? $signed(_T_855_10) : $signed(_GEN_190);
  assign _GEN_192 = 4'hb == _T_659 ? $signed(_T_855_11) : $signed(_GEN_191);
  assign _GEN_193 = 4'hc == _T_659 ? $signed(_T_855_12) : $signed(_GEN_192);
  assign _GEN_194 = 4'hd == _T_659 ? $signed(_T_855_13) : $signed(_GEN_193);
  assign _GEN_195 = 4'he == _T_659 ? $signed(_T_855_14) : $signed(_GEN_194);
  assign _GEN_196 = 4'hf == _T_659 ? $signed(_T_855_15) : $signed(_GEN_195);
  assign _GEN_11 = _GEN_211;
  assign _GEN_197 = 4'h1 == _T_660 ? $signed(_T_925_1) : $signed(_T_925_0);
  assign _GEN_198 = 4'h2 == _T_660 ? $signed(_T_925_2) : $signed(_GEN_197);
  assign _GEN_199 = 4'h3 == _T_660 ? $signed(_T_925_3) : $signed(_GEN_198);
  assign _GEN_200 = 4'h4 == _T_660 ? $signed(_T_925_4) : $signed(_GEN_199);
  assign _GEN_201 = 4'h5 == _T_660 ? $signed(_T_925_5) : $signed(_GEN_200);
  assign _GEN_202 = 4'h6 == _T_660 ? $signed(_T_925_6) : $signed(_GEN_201);
  assign _GEN_203 = 4'h7 == _T_660 ? $signed(_T_925_7) : $signed(_GEN_202);
  assign _GEN_204 = 4'h8 == _T_660 ? $signed(_T_925_8) : $signed(_GEN_203);
  assign _GEN_205 = 4'h9 == _T_660 ? $signed(_T_925_9) : $signed(_GEN_204);
  assign _GEN_206 = 4'ha == _T_660 ? $signed(_T_925_10) : $signed(_GEN_205);
  assign _GEN_207 = 4'hb == _T_660 ? $signed(_T_925_11) : $signed(_GEN_206);
  assign _GEN_208 = 4'hc == _T_660 ? $signed(_T_925_12) : $signed(_GEN_207);
  assign _GEN_209 = 4'hd == _T_660 ? $signed(_T_925_13) : $signed(_GEN_208);
  assign _GEN_210 = 4'he == _T_660 ? $signed(_T_925_14) : $signed(_GEN_209);
  assign _GEN_211 = 4'hf == _T_660 ? $signed(_T_925_15) : $signed(_GEN_210);
  assign _T_1228 = $signed(_GEN_10) + $signed(_GEN_11);
  assign _T_1229 = _T_1228[5:0];
  assign _T_1230 = $signed(_T_1229);
  assign _GEN_12 = _GEN_226;
  assign _GEN_212 = 4'h1 == _T_661 ? $signed(_T_995_1) : $signed(_T_995_0);
  assign _GEN_213 = 4'h2 == _T_661 ? $signed(_T_995_2) : $signed(_GEN_212);
  assign _GEN_214 = 4'h3 == _T_661 ? $signed(_T_995_3) : $signed(_GEN_213);
  assign _GEN_215 = 4'h4 == _T_661 ? $signed(_T_995_4) : $signed(_GEN_214);
  assign _GEN_216 = 4'h5 == _T_661 ? $signed(_T_995_5) : $signed(_GEN_215);
  assign _GEN_217 = 4'h6 == _T_661 ? $signed(_T_995_6) : $signed(_GEN_216);
  assign _GEN_218 = 4'h7 == _T_661 ? $signed(_T_995_7) : $signed(_GEN_217);
  assign _GEN_219 = 4'h8 == _T_661 ? $signed(_T_995_8) : $signed(_GEN_218);
  assign _GEN_220 = 4'h9 == _T_661 ? $signed(_T_995_9) : $signed(_GEN_219);
  assign _GEN_221 = 4'ha == _T_661 ? $signed(_T_995_10) : $signed(_GEN_220);
  assign _GEN_222 = 4'hb == _T_661 ? $signed(_T_995_11) : $signed(_GEN_221);
  assign _GEN_223 = 4'hc == _T_661 ? $signed(_T_995_12) : $signed(_GEN_222);
  assign _GEN_224 = 4'hd == _T_661 ? $signed(_T_995_13) : $signed(_GEN_223);
  assign _GEN_225 = 4'he == _T_661 ? $signed(_T_995_14) : $signed(_GEN_224);
  assign _GEN_226 = 4'hf == _T_661 ? $signed(_T_995_15) : $signed(_GEN_225);
  assign _GEN_13 = _GEN_241;
  assign _GEN_227 = 4'h1 == _T_662 ? $signed(_T_1065_1) : $signed(_T_1065_0);
  assign _GEN_228 = 4'h2 == _T_662 ? $signed(_T_1065_2) : $signed(_GEN_227);
  assign _GEN_229 = 4'h3 == _T_662 ? $signed(_T_1065_3) : $signed(_GEN_228);
  assign _GEN_230 = 4'h4 == _T_662 ? $signed(_T_1065_4) : $signed(_GEN_229);
  assign _GEN_231 = 4'h5 == _T_662 ? $signed(_T_1065_5) : $signed(_GEN_230);
  assign _GEN_232 = 4'h6 == _T_662 ? $signed(_T_1065_6) : $signed(_GEN_231);
  assign _GEN_233 = 4'h7 == _T_662 ? $signed(_T_1065_7) : $signed(_GEN_232);
  assign _GEN_234 = 4'h8 == _T_662 ? $signed(_T_1065_8) : $signed(_GEN_233);
  assign _GEN_235 = 4'h9 == _T_662 ? $signed(_T_1065_9) : $signed(_GEN_234);
  assign _GEN_236 = 4'ha == _T_662 ? $signed(_T_1065_10) : $signed(_GEN_235);
  assign _GEN_237 = 4'hb == _T_662 ? $signed(_T_1065_11) : $signed(_GEN_236);
  assign _GEN_238 = 4'hc == _T_662 ? $signed(_T_1065_12) : $signed(_GEN_237);
  assign _GEN_239 = 4'hd == _T_662 ? $signed(_T_1065_13) : $signed(_GEN_238);
  assign _GEN_240 = 4'he == _T_662 ? $signed(_T_1065_14) : $signed(_GEN_239);
  assign _GEN_241 = 4'hf == _T_662 ? $signed(_T_1065_15) : $signed(_GEN_240);
  assign _T_1231 = $signed(_GEN_12) + $signed(_GEN_13);
  assign _T_1232 = _T_1231[5:0];
  assign _T_1233 = $signed(_T_1232);
  assign _GEN_14 = _GEN_256;
  assign _GEN_242 = 4'h1 == _T_663 ? $signed(_T_1135_1) : $signed(_T_1135_0);
  assign _GEN_243 = 4'h2 == _T_663 ? $signed(_T_1135_2) : $signed(_GEN_242);
  assign _GEN_244 = 4'h3 == _T_663 ? $signed(_T_1135_3) : $signed(_GEN_243);
  assign _GEN_245 = 4'h4 == _T_663 ? $signed(_T_1135_4) : $signed(_GEN_244);
  assign _GEN_246 = 4'h5 == _T_663 ? $signed(_T_1135_5) : $signed(_GEN_245);
  assign _GEN_247 = 4'h6 == _T_663 ? $signed(_T_1135_6) : $signed(_GEN_246);
  assign _GEN_248 = 4'h7 == _T_663 ? $signed(_T_1135_7) : $signed(_GEN_247);
  assign _GEN_249 = 4'h8 == _T_663 ? $signed(_T_1135_8) : $signed(_GEN_248);
  assign _GEN_250 = 4'h9 == _T_663 ? $signed(_T_1135_9) : $signed(_GEN_249);
  assign _GEN_251 = 4'ha == _T_663 ? $signed(_T_1135_10) : $signed(_GEN_250);
  assign _GEN_252 = 4'hb == _T_663 ? $signed(_T_1135_11) : $signed(_GEN_251);
  assign _GEN_253 = 4'hc == _T_663 ? $signed(_T_1135_12) : $signed(_GEN_252);
  assign _GEN_254 = 4'hd == _T_663 ? $signed(_T_1135_13) : $signed(_GEN_253);
  assign _GEN_255 = 4'he == _T_663 ? $signed(_T_1135_14) : $signed(_GEN_254);
  assign _GEN_256 = 4'hf == _T_663 ? $signed(_T_1135_15) : $signed(_GEN_255);
  assign _GEN_15 = _GEN_271;
  assign _GEN_257 = 4'h1 == _T_664 ? $signed(_T_1205_1) : $signed(_T_1205_0);
  assign _GEN_258 = 4'h2 == _T_664 ? $signed(_T_1205_2) : $signed(_GEN_257);
  assign _GEN_259 = 4'h3 == _T_664 ? $signed(_T_1205_3) : $signed(_GEN_258);
  assign _GEN_260 = 4'h4 == _T_664 ? $signed(_T_1205_4) : $signed(_GEN_259);
  assign _GEN_261 = 4'h5 == _T_664 ? $signed(_T_1205_5) : $signed(_GEN_260);
  assign _GEN_262 = 4'h6 == _T_664 ? $signed(_T_1205_6) : $signed(_GEN_261);
  assign _GEN_263 = 4'h7 == _T_664 ? $signed(_T_1205_7) : $signed(_GEN_262);
  assign _GEN_264 = 4'h8 == _T_664 ? $signed(_T_1205_8) : $signed(_GEN_263);
  assign _GEN_265 = 4'h9 == _T_664 ? $signed(_T_1205_9) : $signed(_GEN_264);
  assign _GEN_266 = 4'ha == _T_664 ? $signed(_T_1205_10) : $signed(_GEN_265);
  assign _GEN_267 = 4'hb == _T_664 ? $signed(_T_1205_11) : $signed(_GEN_266);
  assign _GEN_268 = 4'hc == _T_664 ? $signed(_T_1205_12) : $signed(_GEN_267);
  assign _GEN_269 = 4'hd == _T_664 ? $signed(_T_1205_13) : $signed(_GEN_268);
  assign _GEN_270 = 4'he == _T_664 ? $signed(_T_1205_14) : $signed(_GEN_269);
  assign _GEN_271 = 4'hf == _T_664 ? $signed(_T_1205_15) : $signed(_GEN_270);
  assign _T_1234 = $signed(_GEN_14) + $signed(_GEN_15);
  assign _T_1235 = _T_1234[5:0];
  assign _T_1236 = $signed(_T_1235);
  assign _T_1237 = $signed(_T_1227) + $signed(_T_1230);
  assign _T_1238 = _T_1237[5:0];
  assign _T_1239 = $signed(_T_1238);
  assign _T_1240 = $signed(_T_1233) + $signed(_T_1236);
  assign _T_1241 = _T_1240[5:0];
  assign _T_1242 = $signed(_T_1241);
  assign _T_1243 = $signed(_T_1239) + $signed(_T_1242);
  assign _T_1244 = _T_1243[5:0];
  assign _T_1245 = $signed(_T_1244);
  assign MulAdd_1_io_a = _T_1248;
  assign MulAdd_1_io_b = Accumulator_1_io_out;
  assign MulAdd_1_io_m = mean_io_output;
  assign MulAdd_1_io_c = _T_1250;
  assign _T_1246 = mem_io_out[95:64];
  assign _T_1247 = _T_1246[31:16];
  assign _T_1248 = $signed(_T_1247);
  assign _T_1249 = _T_1246[15:0];
  assign _T_1250 = $signed(_T_1249);
  assign _T_1251 = MulAdd_1_io_r[31];
  assign signs_1 = ~ _T_1251;
  assign Accumulator_2_clock = clock;
  assign Accumulator_2_reset = reset;
  assign Accumulator_2_io_in = {{4{_T_1840[5]}},_T_1840};
  assign Accumulator_2_io_sel = io_accSel;
  assign Accumulator_2_io_en = io_accEn;
  assign Accumulator_2_io_reset = io_accReset;
  assign _T_1252 = xnor$_io_out_1[3:0];
  assign _T_1253 = xnor$_io_out_1[7:4];
  assign _T_1254 = xnor$_io_out_1[11:8];
  assign _T_1255 = xnor$_io_out_1[15:12];
  assign _T_1256 = xnor$_io_out_1[19:16];
  assign _T_1257 = xnor$_io_out_1[23:20];
  assign _T_1258 = xnor$_io_out_1[27:24];
  assign _T_1259 = xnor$_io_out_1[31:28];
  assign _T_1310_0 = _T_1262;
  assign _T_1310_1 = _T_1265;
  assign _T_1310_2 = _T_1268;
  assign _T_1310_3 = _T_1271;
  assign _T_1310_4 = _T_1274;
  assign _T_1310_5 = _T_1277;
  assign _T_1310_6 = _T_1280;
  assign _T_1310_7 = _T_1283;
  assign _T_1310_8 = _T_1286;
  assign _T_1310_9 = _T_1289;
  assign _T_1310_10 = _T_1292;
  assign _T_1310_11 = _T_1295;
  assign _T_1310_12 = _T_1298;
  assign _T_1310_13 = _T_1301;
  assign _T_1310_14 = _T_1304;
  assign _T_1310_15 = _T_1307;
  assign _T_1380_0 = _T_1332;
  assign _T_1380_1 = _T_1335;
  assign _T_1380_2 = _T_1338;
  assign _T_1380_3 = _T_1341;
  assign _T_1380_4 = _T_1344;
  assign _T_1380_5 = _T_1347;
  assign _T_1380_6 = _T_1350;
  assign _T_1380_7 = _T_1353;
  assign _T_1380_8 = _T_1356;
  assign _T_1380_9 = _T_1359;
  assign _T_1380_10 = _T_1362;
  assign _T_1380_11 = _T_1365;
  assign _T_1380_12 = _T_1368;
  assign _T_1380_13 = _T_1371;
  assign _T_1380_14 = _T_1374;
  assign _T_1380_15 = _T_1377;
  assign _T_1450_0 = _T_1402;
  assign _T_1450_1 = _T_1405;
  assign _T_1450_2 = _T_1408;
  assign _T_1450_3 = _T_1411;
  assign _T_1450_4 = _T_1414;
  assign _T_1450_5 = _T_1417;
  assign _T_1450_6 = _T_1420;
  assign _T_1450_7 = _T_1423;
  assign _T_1450_8 = _T_1426;
  assign _T_1450_9 = _T_1429;
  assign _T_1450_10 = _T_1432;
  assign _T_1450_11 = _T_1435;
  assign _T_1450_12 = _T_1438;
  assign _T_1450_13 = _T_1441;
  assign _T_1450_14 = _T_1444;
  assign _T_1450_15 = _T_1447;
  assign _T_1520_0 = _T_1472;
  assign _T_1520_1 = _T_1475;
  assign _T_1520_2 = _T_1478;
  assign _T_1520_3 = _T_1481;
  assign _T_1520_4 = _T_1484;
  assign _T_1520_5 = _T_1487;
  assign _T_1520_6 = _T_1490;
  assign _T_1520_7 = _T_1493;
  assign _T_1520_8 = _T_1496;
  assign _T_1520_9 = _T_1499;
  assign _T_1520_10 = _T_1502;
  assign _T_1520_11 = _T_1505;
  assign _T_1520_12 = _T_1508;
  assign _T_1520_13 = _T_1511;
  assign _T_1520_14 = _T_1514;
  assign _T_1520_15 = _T_1517;
  assign _T_1590_0 = _T_1542;
  assign _T_1590_1 = _T_1545;
  assign _T_1590_2 = _T_1548;
  assign _T_1590_3 = _T_1551;
  assign _T_1590_4 = _T_1554;
  assign _T_1590_5 = _T_1557;
  assign _T_1590_6 = _T_1560;
  assign _T_1590_7 = _T_1563;
  assign _T_1590_8 = _T_1566;
  assign _T_1590_9 = _T_1569;
  assign _T_1590_10 = _T_1572;
  assign _T_1590_11 = _T_1575;
  assign _T_1590_12 = _T_1578;
  assign _T_1590_13 = _T_1581;
  assign _T_1590_14 = _T_1584;
  assign _T_1590_15 = _T_1587;
  assign _T_1660_0 = _T_1612;
  assign _T_1660_1 = _T_1615;
  assign _T_1660_2 = _T_1618;
  assign _T_1660_3 = _T_1621;
  assign _T_1660_4 = _T_1624;
  assign _T_1660_5 = _T_1627;
  assign _T_1660_6 = _T_1630;
  assign _T_1660_7 = _T_1633;
  assign _T_1660_8 = _T_1636;
  assign _T_1660_9 = _T_1639;
  assign _T_1660_10 = _T_1642;
  assign _T_1660_11 = _T_1645;
  assign _T_1660_12 = _T_1648;
  assign _T_1660_13 = _T_1651;
  assign _T_1660_14 = _T_1654;
  assign _T_1660_15 = _T_1657;
  assign _T_1730_0 = _T_1682;
  assign _T_1730_1 = _T_1685;
  assign _T_1730_2 = _T_1688;
  assign _T_1730_3 = _T_1691;
  assign _T_1730_4 = _T_1694;
  assign _T_1730_5 = _T_1697;
  assign _T_1730_6 = _T_1700;
  assign _T_1730_7 = _T_1703;
  assign _T_1730_8 = _T_1706;
  assign _T_1730_9 = _T_1709;
  assign _T_1730_10 = _T_1712;
  assign _T_1730_11 = _T_1715;
  assign _T_1730_12 = _T_1718;
  assign _T_1730_13 = _T_1721;
  assign _T_1730_14 = _T_1724;
  assign _T_1730_15 = _T_1727;
  assign _T_1800_0 = _T_1752;
  assign _T_1800_1 = _T_1755;
  assign _T_1800_2 = _T_1758;
  assign _T_1800_3 = _T_1761;
  assign _T_1800_4 = _T_1764;
  assign _T_1800_5 = _T_1767;
  assign _T_1800_6 = _T_1770;
  assign _T_1800_7 = _T_1773;
  assign _T_1800_8 = _T_1776;
  assign _T_1800_9 = _T_1779;
  assign _T_1800_10 = _T_1782;
  assign _T_1800_11 = _T_1785;
  assign _T_1800_12 = _T_1788;
  assign _T_1800_13 = _T_1791;
  assign _T_1800_14 = _T_1794;
  assign _T_1800_15 = _T_1797;
  assign _GEN_16 = _GEN_286;
  assign _GEN_272 = 4'h1 == _T_1252 ? $signed(_T_1310_1) : $signed(_T_1310_0);
  assign _GEN_273 = 4'h2 == _T_1252 ? $signed(_T_1310_2) : $signed(_GEN_272);
  assign _GEN_274 = 4'h3 == _T_1252 ? $signed(_T_1310_3) : $signed(_GEN_273);
  assign _GEN_275 = 4'h4 == _T_1252 ? $signed(_T_1310_4) : $signed(_GEN_274);
  assign _GEN_276 = 4'h5 == _T_1252 ? $signed(_T_1310_5) : $signed(_GEN_275);
  assign _GEN_277 = 4'h6 == _T_1252 ? $signed(_T_1310_6) : $signed(_GEN_276);
  assign _GEN_278 = 4'h7 == _T_1252 ? $signed(_T_1310_7) : $signed(_GEN_277);
  assign _GEN_279 = 4'h8 == _T_1252 ? $signed(_T_1310_8) : $signed(_GEN_278);
  assign _GEN_280 = 4'h9 == _T_1252 ? $signed(_T_1310_9) : $signed(_GEN_279);
  assign _GEN_281 = 4'ha == _T_1252 ? $signed(_T_1310_10) : $signed(_GEN_280);
  assign _GEN_282 = 4'hb == _T_1252 ? $signed(_T_1310_11) : $signed(_GEN_281);
  assign _GEN_283 = 4'hc == _T_1252 ? $signed(_T_1310_12) : $signed(_GEN_282);
  assign _GEN_284 = 4'hd == _T_1252 ? $signed(_T_1310_13) : $signed(_GEN_283);
  assign _GEN_285 = 4'he == _T_1252 ? $signed(_T_1310_14) : $signed(_GEN_284);
  assign _GEN_286 = 4'hf == _T_1252 ? $signed(_T_1310_15) : $signed(_GEN_285);
  assign _GEN_17 = _GEN_301;
  assign _GEN_287 = 4'h1 == _T_1253 ? $signed(_T_1380_1) : $signed(_T_1380_0);
  assign _GEN_288 = 4'h2 == _T_1253 ? $signed(_T_1380_2) : $signed(_GEN_287);
  assign _GEN_289 = 4'h3 == _T_1253 ? $signed(_T_1380_3) : $signed(_GEN_288);
  assign _GEN_290 = 4'h4 == _T_1253 ? $signed(_T_1380_4) : $signed(_GEN_289);
  assign _GEN_291 = 4'h5 == _T_1253 ? $signed(_T_1380_5) : $signed(_GEN_290);
  assign _GEN_292 = 4'h6 == _T_1253 ? $signed(_T_1380_6) : $signed(_GEN_291);
  assign _GEN_293 = 4'h7 == _T_1253 ? $signed(_T_1380_7) : $signed(_GEN_292);
  assign _GEN_294 = 4'h8 == _T_1253 ? $signed(_T_1380_8) : $signed(_GEN_293);
  assign _GEN_295 = 4'h9 == _T_1253 ? $signed(_T_1380_9) : $signed(_GEN_294);
  assign _GEN_296 = 4'ha == _T_1253 ? $signed(_T_1380_10) : $signed(_GEN_295);
  assign _GEN_297 = 4'hb == _T_1253 ? $signed(_T_1380_11) : $signed(_GEN_296);
  assign _GEN_298 = 4'hc == _T_1253 ? $signed(_T_1380_12) : $signed(_GEN_297);
  assign _GEN_299 = 4'hd == _T_1253 ? $signed(_T_1380_13) : $signed(_GEN_298);
  assign _GEN_300 = 4'he == _T_1253 ? $signed(_T_1380_14) : $signed(_GEN_299);
  assign _GEN_301 = 4'hf == _T_1253 ? $signed(_T_1380_15) : $signed(_GEN_300);
  assign _T_1820 = $signed(_GEN_16) + $signed(_GEN_17);
  assign _T_1821 = _T_1820[5:0];
  assign _T_1822 = $signed(_T_1821);
  assign _GEN_18 = _GEN_316;
  assign _GEN_302 = 4'h1 == _T_1254 ? $signed(_T_1450_1) : $signed(_T_1450_0);
  assign _GEN_303 = 4'h2 == _T_1254 ? $signed(_T_1450_2) : $signed(_GEN_302);
  assign _GEN_304 = 4'h3 == _T_1254 ? $signed(_T_1450_3) : $signed(_GEN_303);
  assign _GEN_305 = 4'h4 == _T_1254 ? $signed(_T_1450_4) : $signed(_GEN_304);
  assign _GEN_306 = 4'h5 == _T_1254 ? $signed(_T_1450_5) : $signed(_GEN_305);
  assign _GEN_307 = 4'h6 == _T_1254 ? $signed(_T_1450_6) : $signed(_GEN_306);
  assign _GEN_308 = 4'h7 == _T_1254 ? $signed(_T_1450_7) : $signed(_GEN_307);
  assign _GEN_309 = 4'h8 == _T_1254 ? $signed(_T_1450_8) : $signed(_GEN_308);
  assign _GEN_310 = 4'h9 == _T_1254 ? $signed(_T_1450_9) : $signed(_GEN_309);
  assign _GEN_311 = 4'ha == _T_1254 ? $signed(_T_1450_10) : $signed(_GEN_310);
  assign _GEN_312 = 4'hb == _T_1254 ? $signed(_T_1450_11) : $signed(_GEN_311);
  assign _GEN_313 = 4'hc == _T_1254 ? $signed(_T_1450_12) : $signed(_GEN_312);
  assign _GEN_314 = 4'hd == _T_1254 ? $signed(_T_1450_13) : $signed(_GEN_313);
  assign _GEN_315 = 4'he == _T_1254 ? $signed(_T_1450_14) : $signed(_GEN_314);
  assign _GEN_316 = 4'hf == _T_1254 ? $signed(_T_1450_15) : $signed(_GEN_315);
  assign _GEN_19 = _GEN_331;
  assign _GEN_317 = 4'h1 == _T_1255 ? $signed(_T_1520_1) : $signed(_T_1520_0);
  assign _GEN_318 = 4'h2 == _T_1255 ? $signed(_T_1520_2) : $signed(_GEN_317);
  assign _GEN_319 = 4'h3 == _T_1255 ? $signed(_T_1520_3) : $signed(_GEN_318);
  assign _GEN_320 = 4'h4 == _T_1255 ? $signed(_T_1520_4) : $signed(_GEN_319);
  assign _GEN_321 = 4'h5 == _T_1255 ? $signed(_T_1520_5) : $signed(_GEN_320);
  assign _GEN_322 = 4'h6 == _T_1255 ? $signed(_T_1520_6) : $signed(_GEN_321);
  assign _GEN_323 = 4'h7 == _T_1255 ? $signed(_T_1520_7) : $signed(_GEN_322);
  assign _GEN_324 = 4'h8 == _T_1255 ? $signed(_T_1520_8) : $signed(_GEN_323);
  assign _GEN_325 = 4'h9 == _T_1255 ? $signed(_T_1520_9) : $signed(_GEN_324);
  assign _GEN_326 = 4'ha == _T_1255 ? $signed(_T_1520_10) : $signed(_GEN_325);
  assign _GEN_327 = 4'hb == _T_1255 ? $signed(_T_1520_11) : $signed(_GEN_326);
  assign _GEN_328 = 4'hc == _T_1255 ? $signed(_T_1520_12) : $signed(_GEN_327);
  assign _GEN_329 = 4'hd == _T_1255 ? $signed(_T_1520_13) : $signed(_GEN_328);
  assign _GEN_330 = 4'he == _T_1255 ? $signed(_T_1520_14) : $signed(_GEN_329);
  assign _GEN_331 = 4'hf == _T_1255 ? $signed(_T_1520_15) : $signed(_GEN_330);
  assign _T_1823 = $signed(_GEN_18) + $signed(_GEN_19);
  assign _T_1824 = _T_1823[5:0];
  assign _T_1825 = $signed(_T_1824);
  assign _GEN_20 = _GEN_346;
  assign _GEN_332 = 4'h1 == _T_1256 ? $signed(_T_1590_1) : $signed(_T_1590_0);
  assign _GEN_333 = 4'h2 == _T_1256 ? $signed(_T_1590_2) : $signed(_GEN_332);
  assign _GEN_334 = 4'h3 == _T_1256 ? $signed(_T_1590_3) : $signed(_GEN_333);
  assign _GEN_335 = 4'h4 == _T_1256 ? $signed(_T_1590_4) : $signed(_GEN_334);
  assign _GEN_336 = 4'h5 == _T_1256 ? $signed(_T_1590_5) : $signed(_GEN_335);
  assign _GEN_337 = 4'h6 == _T_1256 ? $signed(_T_1590_6) : $signed(_GEN_336);
  assign _GEN_338 = 4'h7 == _T_1256 ? $signed(_T_1590_7) : $signed(_GEN_337);
  assign _GEN_339 = 4'h8 == _T_1256 ? $signed(_T_1590_8) : $signed(_GEN_338);
  assign _GEN_340 = 4'h9 == _T_1256 ? $signed(_T_1590_9) : $signed(_GEN_339);
  assign _GEN_341 = 4'ha == _T_1256 ? $signed(_T_1590_10) : $signed(_GEN_340);
  assign _GEN_342 = 4'hb == _T_1256 ? $signed(_T_1590_11) : $signed(_GEN_341);
  assign _GEN_343 = 4'hc == _T_1256 ? $signed(_T_1590_12) : $signed(_GEN_342);
  assign _GEN_344 = 4'hd == _T_1256 ? $signed(_T_1590_13) : $signed(_GEN_343);
  assign _GEN_345 = 4'he == _T_1256 ? $signed(_T_1590_14) : $signed(_GEN_344);
  assign _GEN_346 = 4'hf == _T_1256 ? $signed(_T_1590_15) : $signed(_GEN_345);
  assign _GEN_21 = _GEN_361;
  assign _GEN_347 = 4'h1 == _T_1257 ? $signed(_T_1660_1) : $signed(_T_1660_0);
  assign _GEN_348 = 4'h2 == _T_1257 ? $signed(_T_1660_2) : $signed(_GEN_347);
  assign _GEN_349 = 4'h3 == _T_1257 ? $signed(_T_1660_3) : $signed(_GEN_348);
  assign _GEN_350 = 4'h4 == _T_1257 ? $signed(_T_1660_4) : $signed(_GEN_349);
  assign _GEN_351 = 4'h5 == _T_1257 ? $signed(_T_1660_5) : $signed(_GEN_350);
  assign _GEN_352 = 4'h6 == _T_1257 ? $signed(_T_1660_6) : $signed(_GEN_351);
  assign _GEN_353 = 4'h7 == _T_1257 ? $signed(_T_1660_7) : $signed(_GEN_352);
  assign _GEN_354 = 4'h8 == _T_1257 ? $signed(_T_1660_8) : $signed(_GEN_353);
  assign _GEN_355 = 4'h9 == _T_1257 ? $signed(_T_1660_9) : $signed(_GEN_354);
  assign _GEN_356 = 4'ha == _T_1257 ? $signed(_T_1660_10) : $signed(_GEN_355);
  assign _GEN_357 = 4'hb == _T_1257 ? $signed(_T_1660_11) : $signed(_GEN_356);
  assign _GEN_358 = 4'hc == _T_1257 ? $signed(_T_1660_12) : $signed(_GEN_357);
  assign _GEN_359 = 4'hd == _T_1257 ? $signed(_T_1660_13) : $signed(_GEN_358);
  assign _GEN_360 = 4'he == _T_1257 ? $signed(_T_1660_14) : $signed(_GEN_359);
  assign _GEN_361 = 4'hf == _T_1257 ? $signed(_T_1660_15) : $signed(_GEN_360);
  assign _T_1826 = $signed(_GEN_20) + $signed(_GEN_21);
  assign _T_1827 = _T_1826[5:0];
  assign _T_1828 = $signed(_T_1827);
  assign _GEN_22 = _GEN_376;
  assign _GEN_362 = 4'h1 == _T_1258 ? $signed(_T_1730_1) : $signed(_T_1730_0);
  assign _GEN_363 = 4'h2 == _T_1258 ? $signed(_T_1730_2) : $signed(_GEN_362);
  assign _GEN_364 = 4'h3 == _T_1258 ? $signed(_T_1730_3) : $signed(_GEN_363);
  assign _GEN_365 = 4'h4 == _T_1258 ? $signed(_T_1730_4) : $signed(_GEN_364);
  assign _GEN_366 = 4'h5 == _T_1258 ? $signed(_T_1730_5) : $signed(_GEN_365);
  assign _GEN_367 = 4'h6 == _T_1258 ? $signed(_T_1730_6) : $signed(_GEN_366);
  assign _GEN_368 = 4'h7 == _T_1258 ? $signed(_T_1730_7) : $signed(_GEN_367);
  assign _GEN_369 = 4'h8 == _T_1258 ? $signed(_T_1730_8) : $signed(_GEN_368);
  assign _GEN_370 = 4'h9 == _T_1258 ? $signed(_T_1730_9) : $signed(_GEN_369);
  assign _GEN_371 = 4'ha == _T_1258 ? $signed(_T_1730_10) : $signed(_GEN_370);
  assign _GEN_372 = 4'hb == _T_1258 ? $signed(_T_1730_11) : $signed(_GEN_371);
  assign _GEN_373 = 4'hc == _T_1258 ? $signed(_T_1730_12) : $signed(_GEN_372);
  assign _GEN_374 = 4'hd == _T_1258 ? $signed(_T_1730_13) : $signed(_GEN_373);
  assign _GEN_375 = 4'he == _T_1258 ? $signed(_T_1730_14) : $signed(_GEN_374);
  assign _GEN_376 = 4'hf == _T_1258 ? $signed(_T_1730_15) : $signed(_GEN_375);
  assign _GEN_23 = _GEN_391;
  assign _GEN_377 = 4'h1 == _T_1259 ? $signed(_T_1800_1) : $signed(_T_1800_0);
  assign _GEN_378 = 4'h2 == _T_1259 ? $signed(_T_1800_2) : $signed(_GEN_377);
  assign _GEN_379 = 4'h3 == _T_1259 ? $signed(_T_1800_3) : $signed(_GEN_378);
  assign _GEN_380 = 4'h4 == _T_1259 ? $signed(_T_1800_4) : $signed(_GEN_379);
  assign _GEN_381 = 4'h5 == _T_1259 ? $signed(_T_1800_5) : $signed(_GEN_380);
  assign _GEN_382 = 4'h6 == _T_1259 ? $signed(_T_1800_6) : $signed(_GEN_381);
  assign _GEN_383 = 4'h7 == _T_1259 ? $signed(_T_1800_7) : $signed(_GEN_382);
  assign _GEN_384 = 4'h8 == _T_1259 ? $signed(_T_1800_8) : $signed(_GEN_383);
  assign _GEN_385 = 4'h9 == _T_1259 ? $signed(_T_1800_9) : $signed(_GEN_384);
  assign _GEN_386 = 4'ha == _T_1259 ? $signed(_T_1800_10) : $signed(_GEN_385);
  assign _GEN_387 = 4'hb == _T_1259 ? $signed(_T_1800_11) : $signed(_GEN_386);
  assign _GEN_388 = 4'hc == _T_1259 ? $signed(_T_1800_12) : $signed(_GEN_387);
  assign _GEN_389 = 4'hd == _T_1259 ? $signed(_T_1800_13) : $signed(_GEN_388);
  assign _GEN_390 = 4'he == _T_1259 ? $signed(_T_1800_14) : $signed(_GEN_389);
  assign _GEN_391 = 4'hf == _T_1259 ? $signed(_T_1800_15) : $signed(_GEN_390);
  assign _T_1829 = $signed(_GEN_22) + $signed(_GEN_23);
  assign _T_1830 = _T_1829[5:0];
  assign _T_1831 = $signed(_T_1830);
  assign _T_1832 = $signed(_T_1822) + $signed(_T_1825);
  assign _T_1833 = _T_1832[5:0];
  assign _T_1834 = $signed(_T_1833);
  assign _T_1835 = $signed(_T_1828) + $signed(_T_1831);
  assign _T_1836 = _T_1835[5:0];
  assign _T_1837 = $signed(_T_1836);
  assign _T_1838 = $signed(_T_1834) + $signed(_T_1837);
  assign _T_1839 = _T_1838[5:0];
  assign _T_1840 = $signed(_T_1839);
  assign MulAdd_2_io_a = _T_1843;
  assign MulAdd_2_io_b = Accumulator_2_io_out;
  assign MulAdd_2_io_m = mean_io_output;
  assign MulAdd_2_io_c = _T_1845;
  assign _T_1841 = mem_io_out[63:32];
  assign _T_1842 = _T_1841[31:16];
  assign _T_1843 = $signed(_T_1842);
  assign _T_1844 = _T_1841[15:0];
  assign _T_1845 = $signed(_T_1844);
  assign _T_1846 = MulAdd_2_io_r[31];
  assign signs_2 = ~ _T_1846;
  assign Accumulator_3_clock = clock;
  assign Accumulator_3_reset = reset;
  assign Accumulator_3_io_in = {{4{_T_2435[5]}},_T_2435};
  assign Accumulator_3_io_sel = io_accSel;
  assign Accumulator_3_io_en = io_accEn;
  assign Accumulator_3_io_reset = io_accReset;
  assign _T_1847 = xnor$_io_out_0[3:0];
  assign _T_1848 = xnor$_io_out_0[7:4];
  assign _T_1849 = xnor$_io_out_0[11:8];
  assign _T_1850 = xnor$_io_out_0[15:12];
  assign _T_1851 = xnor$_io_out_0[19:16];
  assign _T_1852 = xnor$_io_out_0[23:20];
  assign _T_1853 = xnor$_io_out_0[27:24];
  assign _T_1854 = xnor$_io_out_0[31:28];
  assign _T_1905_0 = _T_1857;
  assign _T_1905_1 = _T_1860;
  assign _T_1905_2 = _T_1863;
  assign _T_1905_3 = _T_1866;
  assign _T_1905_4 = _T_1869;
  assign _T_1905_5 = _T_1872;
  assign _T_1905_6 = _T_1875;
  assign _T_1905_7 = _T_1878;
  assign _T_1905_8 = _T_1881;
  assign _T_1905_9 = _T_1884;
  assign _T_1905_10 = _T_1887;
  assign _T_1905_11 = _T_1890;
  assign _T_1905_12 = _T_1893;
  assign _T_1905_13 = _T_1896;
  assign _T_1905_14 = _T_1899;
  assign _T_1905_15 = _T_1902;
  assign _T_1975_0 = _T_1927;
  assign _T_1975_1 = _T_1930;
  assign _T_1975_2 = _T_1933;
  assign _T_1975_3 = _T_1936;
  assign _T_1975_4 = _T_1939;
  assign _T_1975_5 = _T_1942;
  assign _T_1975_6 = _T_1945;
  assign _T_1975_7 = _T_1948;
  assign _T_1975_8 = _T_1951;
  assign _T_1975_9 = _T_1954;
  assign _T_1975_10 = _T_1957;
  assign _T_1975_11 = _T_1960;
  assign _T_1975_12 = _T_1963;
  assign _T_1975_13 = _T_1966;
  assign _T_1975_14 = _T_1969;
  assign _T_1975_15 = _T_1972;
  assign _T_2045_0 = _T_1997;
  assign _T_2045_1 = _T_2000;
  assign _T_2045_2 = _T_2003;
  assign _T_2045_3 = _T_2006;
  assign _T_2045_4 = _T_2009;
  assign _T_2045_5 = _T_2012;
  assign _T_2045_6 = _T_2015;
  assign _T_2045_7 = _T_2018;
  assign _T_2045_8 = _T_2021;
  assign _T_2045_9 = _T_2024;
  assign _T_2045_10 = _T_2027;
  assign _T_2045_11 = _T_2030;
  assign _T_2045_12 = _T_2033;
  assign _T_2045_13 = _T_2036;
  assign _T_2045_14 = _T_2039;
  assign _T_2045_15 = _T_2042;
  assign _T_2115_0 = _T_2067;
  assign _T_2115_1 = _T_2070;
  assign _T_2115_2 = _T_2073;
  assign _T_2115_3 = _T_2076;
  assign _T_2115_4 = _T_2079;
  assign _T_2115_5 = _T_2082;
  assign _T_2115_6 = _T_2085;
  assign _T_2115_7 = _T_2088;
  assign _T_2115_8 = _T_2091;
  assign _T_2115_9 = _T_2094;
  assign _T_2115_10 = _T_2097;
  assign _T_2115_11 = _T_2100;
  assign _T_2115_12 = _T_2103;
  assign _T_2115_13 = _T_2106;
  assign _T_2115_14 = _T_2109;
  assign _T_2115_15 = _T_2112;
  assign _T_2185_0 = _T_2137;
  assign _T_2185_1 = _T_2140;
  assign _T_2185_2 = _T_2143;
  assign _T_2185_3 = _T_2146;
  assign _T_2185_4 = _T_2149;
  assign _T_2185_5 = _T_2152;
  assign _T_2185_6 = _T_2155;
  assign _T_2185_7 = _T_2158;
  assign _T_2185_8 = _T_2161;
  assign _T_2185_9 = _T_2164;
  assign _T_2185_10 = _T_2167;
  assign _T_2185_11 = _T_2170;
  assign _T_2185_12 = _T_2173;
  assign _T_2185_13 = _T_2176;
  assign _T_2185_14 = _T_2179;
  assign _T_2185_15 = _T_2182;
  assign _T_2255_0 = _T_2207;
  assign _T_2255_1 = _T_2210;
  assign _T_2255_2 = _T_2213;
  assign _T_2255_3 = _T_2216;
  assign _T_2255_4 = _T_2219;
  assign _T_2255_5 = _T_2222;
  assign _T_2255_6 = _T_2225;
  assign _T_2255_7 = _T_2228;
  assign _T_2255_8 = _T_2231;
  assign _T_2255_9 = _T_2234;
  assign _T_2255_10 = _T_2237;
  assign _T_2255_11 = _T_2240;
  assign _T_2255_12 = _T_2243;
  assign _T_2255_13 = _T_2246;
  assign _T_2255_14 = _T_2249;
  assign _T_2255_15 = _T_2252;
  assign _T_2325_0 = _T_2277;
  assign _T_2325_1 = _T_2280;
  assign _T_2325_2 = _T_2283;
  assign _T_2325_3 = _T_2286;
  assign _T_2325_4 = _T_2289;
  assign _T_2325_5 = _T_2292;
  assign _T_2325_6 = _T_2295;
  assign _T_2325_7 = _T_2298;
  assign _T_2325_8 = _T_2301;
  assign _T_2325_9 = _T_2304;
  assign _T_2325_10 = _T_2307;
  assign _T_2325_11 = _T_2310;
  assign _T_2325_12 = _T_2313;
  assign _T_2325_13 = _T_2316;
  assign _T_2325_14 = _T_2319;
  assign _T_2325_15 = _T_2322;
  assign _T_2395_0 = _T_2347;
  assign _T_2395_1 = _T_2350;
  assign _T_2395_2 = _T_2353;
  assign _T_2395_3 = _T_2356;
  assign _T_2395_4 = _T_2359;
  assign _T_2395_5 = _T_2362;
  assign _T_2395_6 = _T_2365;
  assign _T_2395_7 = _T_2368;
  assign _T_2395_8 = _T_2371;
  assign _T_2395_9 = _T_2374;
  assign _T_2395_10 = _T_2377;
  assign _T_2395_11 = _T_2380;
  assign _T_2395_12 = _T_2383;
  assign _T_2395_13 = _T_2386;
  assign _T_2395_14 = _T_2389;
  assign _T_2395_15 = _T_2392;
  assign _GEN_24 = _GEN_406;
  assign _GEN_392 = 4'h1 == _T_1847 ? $signed(_T_1905_1) : $signed(_T_1905_0);
  assign _GEN_393 = 4'h2 == _T_1847 ? $signed(_T_1905_2) : $signed(_GEN_392);
  assign _GEN_394 = 4'h3 == _T_1847 ? $signed(_T_1905_3) : $signed(_GEN_393);
  assign _GEN_395 = 4'h4 == _T_1847 ? $signed(_T_1905_4) : $signed(_GEN_394);
  assign _GEN_396 = 4'h5 == _T_1847 ? $signed(_T_1905_5) : $signed(_GEN_395);
  assign _GEN_397 = 4'h6 == _T_1847 ? $signed(_T_1905_6) : $signed(_GEN_396);
  assign _GEN_398 = 4'h7 == _T_1847 ? $signed(_T_1905_7) : $signed(_GEN_397);
  assign _GEN_399 = 4'h8 == _T_1847 ? $signed(_T_1905_8) : $signed(_GEN_398);
  assign _GEN_400 = 4'h9 == _T_1847 ? $signed(_T_1905_9) : $signed(_GEN_399);
  assign _GEN_401 = 4'ha == _T_1847 ? $signed(_T_1905_10) : $signed(_GEN_400);
  assign _GEN_402 = 4'hb == _T_1847 ? $signed(_T_1905_11) : $signed(_GEN_401);
  assign _GEN_403 = 4'hc == _T_1847 ? $signed(_T_1905_12) : $signed(_GEN_402);
  assign _GEN_404 = 4'hd == _T_1847 ? $signed(_T_1905_13) : $signed(_GEN_403);
  assign _GEN_405 = 4'he == _T_1847 ? $signed(_T_1905_14) : $signed(_GEN_404);
  assign _GEN_406 = 4'hf == _T_1847 ? $signed(_T_1905_15) : $signed(_GEN_405);
  assign _GEN_25 = _GEN_421;
  assign _GEN_407 = 4'h1 == _T_1848 ? $signed(_T_1975_1) : $signed(_T_1975_0);
  assign _GEN_408 = 4'h2 == _T_1848 ? $signed(_T_1975_2) : $signed(_GEN_407);
  assign _GEN_409 = 4'h3 == _T_1848 ? $signed(_T_1975_3) : $signed(_GEN_408);
  assign _GEN_410 = 4'h4 == _T_1848 ? $signed(_T_1975_4) : $signed(_GEN_409);
  assign _GEN_411 = 4'h5 == _T_1848 ? $signed(_T_1975_5) : $signed(_GEN_410);
  assign _GEN_412 = 4'h6 == _T_1848 ? $signed(_T_1975_6) : $signed(_GEN_411);
  assign _GEN_413 = 4'h7 == _T_1848 ? $signed(_T_1975_7) : $signed(_GEN_412);
  assign _GEN_414 = 4'h8 == _T_1848 ? $signed(_T_1975_8) : $signed(_GEN_413);
  assign _GEN_415 = 4'h9 == _T_1848 ? $signed(_T_1975_9) : $signed(_GEN_414);
  assign _GEN_416 = 4'ha == _T_1848 ? $signed(_T_1975_10) : $signed(_GEN_415);
  assign _GEN_417 = 4'hb == _T_1848 ? $signed(_T_1975_11) : $signed(_GEN_416);
  assign _GEN_418 = 4'hc == _T_1848 ? $signed(_T_1975_12) : $signed(_GEN_417);
  assign _GEN_419 = 4'hd == _T_1848 ? $signed(_T_1975_13) : $signed(_GEN_418);
  assign _GEN_420 = 4'he == _T_1848 ? $signed(_T_1975_14) : $signed(_GEN_419);
  assign _GEN_421 = 4'hf == _T_1848 ? $signed(_T_1975_15) : $signed(_GEN_420);
  assign _T_2415 = $signed(_GEN_24) + $signed(_GEN_25);
  assign _T_2416 = _T_2415[5:0];
  assign _T_2417 = $signed(_T_2416);
  assign _GEN_26 = _GEN_436;
  assign _GEN_422 = 4'h1 == _T_1849 ? $signed(_T_2045_1) : $signed(_T_2045_0);
  assign _GEN_423 = 4'h2 == _T_1849 ? $signed(_T_2045_2) : $signed(_GEN_422);
  assign _GEN_424 = 4'h3 == _T_1849 ? $signed(_T_2045_3) : $signed(_GEN_423);
  assign _GEN_425 = 4'h4 == _T_1849 ? $signed(_T_2045_4) : $signed(_GEN_424);
  assign _GEN_426 = 4'h5 == _T_1849 ? $signed(_T_2045_5) : $signed(_GEN_425);
  assign _GEN_427 = 4'h6 == _T_1849 ? $signed(_T_2045_6) : $signed(_GEN_426);
  assign _GEN_428 = 4'h7 == _T_1849 ? $signed(_T_2045_7) : $signed(_GEN_427);
  assign _GEN_429 = 4'h8 == _T_1849 ? $signed(_T_2045_8) : $signed(_GEN_428);
  assign _GEN_430 = 4'h9 == _T_1849 ? $signed(_T_2045_9) : $signed(_GEN_429);
  assign _GEN_431 = 4'ha == _T_1849 ? $signed(_T_2045_10) : $signed(_GEN_430);
  assign _GEN_432 = 4'hb == _T_1849 ? $signed(_T_2045_11) : $signed(_GEN_431);
  assign _GEN_433 = 4'hc == _T_1849 ? $signed(_T_2045_12) : $signed(_GEN_432);
  assign _GEN_434 = 4'hd == _T_1849 ? $signed(_T_2045_13) : $signed(_GEN_433);
  assign _GEN_435 = 4'he == _T_1849 ? $signed(_T_2045_14) : $signed(_GEN_434);
  assign _GEN_436 = 4'hf == _T_1849 ? $signed(_T_2045_15) : $signed(_GEN_435);
  assign _GEN_27 = _GEN_451;
  assign _GEN_437 = 4'h1 == _T_1850 ? $signed(_T_2115_1) : $signed(_T_2115_0);
  assign _GEN_438 = 4'h2 == _T_1850 ? $signed(_T_2115_2) : $signed(_GEN_437);
  assign _GEN_439 = 4'h3 == _T_1850 ? $signed(_T_2115_3) : $signed(_GEN_438);
  assign _GEN_440 = 4'h4 == _T_1850 ? $signed(_T_2115_4) : $signed(_GEN_439);
  assign _GEN_441 = 4'h5 == _T_1850 ? $signed(_T_2115_5) : $signed(_GEN_440);
  assign _GEN_442 = 4'h6 == _T_1850 ? $signed(_T_2115_6) : $signed(_GEN_441);
  assign _GEN_443 = 4'h7 == _T_1850 ? $signed(_T_2115_7) : $signed(_GEN_442);
  assign _GEN_444 = 4'h8 == _T_1850 ? $signed(_T_2115_8) : $signed(_GEN_443);
  assign _GEN_445 = 4'h9 == _T_1850 ? $signed(_T_2115_9) : $signed(_GEN_444);
  assign _GEN_446 = 4'ha == _T_1850 ? $signed(_T_2115_10) : $signed(_GEN_445);
  assign _GEN_447 = 4'hb == _T_1850 ? $signed(_T_2115_11) : $signed(_GEN_446);
  assign _GEN_448 = 4'hc == _T_1850 ? $signed(_T_2115_12) : $signed(_GEN_447);
  assign _GEN_449 = 4'hd == _T_1850 ? $signed(_T_2115_13) : $signed(_GEN_448);
  assign _GEN_450 = 4'he == _T_1850 ? $signed(_T_2115_14) : $signed(_GEN_449);
  assign _GEN_451 = 4'hf == _T_1850 ? $signed(_T_2115_15) : $signed(_GEN_450);
  assign _T_2418 = $signed(_GEN_26) + $signed(_GEN_27);
  assign _T_2419 = _T_2418[5:0];
  assign _T_2420 = $signed(_T_2419);
  assign _GEN_28 = _GEN_466;
  assign _GEN_452 = 4'h1 == _T_1851 ? $signed(_T_2185_1) : $signed(_T_2185_0);
  assign _GEN_453 = 4'h2 == _T_1851 ? $signed(_T_2185_2) : $signed(_GEN_452);
  assign _GEN_454 = 4'h3 == _T_1851 ? $signed(_T_2185_3) : $signed(_GEN_453);
  assign _GEN_455 = 4'h4 == _T_1851 ? $signed(_T_2185_4) : $signed(_GEN_454);
  assign _GEN_456 = 4'h5 == _T_1851 ? $signed(_T_2185_5) : $signed(_GEN_455);
  assign _GEN_457 = 4'h6 == _T_1851 ? $signed(_T_2185_6) : $signed(_GEN_456);
  assign _GEN_458 = 4'h7 == _T_1851 ? $signed(_T_2185_7) : $signed(_GEN_457);
  assign _GEN_459 = 4'h8 == _T_1851 ? $signed(_T_2185_8) : $signed(_GEN_458);
  assign _GEN_460 = 4'h9 == _T_1851 ? $signed(_T_2185_9) : $signed(_GEN_459);
  assign _GEN_461 = 4'ha == _T_1851 ? $signed(_T_2185_10) : $signed(_GEN_460);
  assign _GEN_462 = 4'hb == _T_1851 ? $signed(_T_2185_11) : $signed(_GEN_461);
  assign _GEN_463 = 4'hc == _T_1851 ? $signed(_T_2185_12) : $signed(_GEN_462);
  assign _GEN_464 = 4'hd == _T_1851 ? $signed(_T_2185_13) : $signed(_GEN_463);
  assign _GEN_465 = 4'he == _T_1851 ? $signed(_T_2185_14) : $signed(_GEN_464);
  assign _GEN_466 = 4'hf == _T_1851 ? $signed(_T_2185_15) : $signed(_GEN_465);
  assign _GEN_29 = _GEN_481;
  assign _GEN_467 = 4'h1 == _T_1852 ? $signed(_T_2255_1) : $signed(_T_2255_0);
  assign _GEN_468 = 4'h2 == _T_1852 ? $signed(_T_2255_2) : $signed(_GEN_467);
  assign _GEN_469 = 4'h3 == _T_1852 ? $signed(_T_2255_3) : $signed(_GEN_468);
  assign _GEN_470 = 4'h4 == _T_1852 ? $signed(_T_2255_4) : $signed(_GEN_469);
  assign _GEN_471 = 4'h5 == _T_1852 ? $signed(_T_2255_5) : $signed(_GEN_470);
  assign _GEN_472 = 4'h6 == _T_1852 ? $signed(_T_2255_6) : $signed(_GEN_471);
  assign _GEN_473 = 4'h7 == _T_1852 ? $signed(_T_2255_7) : $signed(_GEN_472);
  assign _GEN_474 = 4'h8 == _T_1852 ? $signed(_T_2255_8) : $signed(_GEN_473);
  assign _GEN_475 = 4'h9 == _T_1852 ? $signed(_T_2255_9) : $signed(_GEN_474);
  assign _GEN_476 = 4'ha == _T_1852 ? $signed(_T_2255_10) : $signed(_GEN_475);
  assign _GEN_477 = 4'hb == _T_1852 ? $signed(_T_2255_11) : $signed(_GEN_476);
  assign _GEN_478 = 4'hc == _T_1852 ? $signed(_T_2255_12) : $signed(_GEN_477);
  assign _GEN_479 = 4'hd == _T_1852 ? $signed(_T_2255_13) : $signed(_GEN_478);
  assign _GEN_480 = 4'he == _T_1852 ? $signed(_T_2255_14) : $signed(_GEN_479);
  assign _GEN_481 = 4'hf == _T_1852 ? $signed(_T_2255_15) : $signed(_GEN_480);
  assign _T_2421 = $signed(_GEN_28) + $signed(_GEN_29);
  assign _T_2422 = _T_2421[5:0];
  assign _T_2423 = $signed(_T_2422);
  assign _GEN_30 = _GEN_496;
  assign _GEN_482 = 4'h1 == _T_1853 ? $signed(_T_2325_1) : $signed(_T_2325_0);
  assign _GEN_483 = 4'h2 == _T_1853 ? $signed(_T_2325_2) : $signed(_GEN_482);
  assign _GEN_484 = 4'h3 == _T_1853 ? $signed(_T_2325_3) : $signed(_GEN_483);
  assign _GEN_485 = 4'h4 == _T_1853 ? $signed(_T_2325_4) : $signed(_GEN_484);
  assign _GEN_486 = 4'h5 == _T_1853 ? $signed(_T_2325_5) : $signed(_GEN_485);
  assign _GEN_487 = 4'h6 == _T_1853 ? $signed(_T_2325_6) : $signed(_GEN_486);
  assign _GEN_488 = 4'h7 == _T_1853 ? $signed(_T_2325_7) : $signed(_GEN_487);
  assign _GEN_489 = 4'h8 == _T_1853 ? $signed(_T_2325_8) : $signed(_GEN_488);
  assign _GEN_490 = 4'h9 == _T_1853 ? $signed(_T_2325_9) : $signed(_GEN_489);
  assign _GEN_491 = 4'ha == _T_1853 ? $signed(_T_2325_10) : $signed(_GEN_490);
  assign _GEN_492 = 4'hb == _T_1853 ? $signed(_T_2325_11) : $signed(_GEN_491);
  assign _GEN_493 = 4'hc == _T_1853 ? $signed(_T_2325_12) : $signed(_GEN_492);
  assign _GEN_494 = 4'hd == _T_1853 ? $signed(_T_2325_13) : $signed(_GEN_493);
  assign _GEN_495 = 4'he == _T_1853 ? $signed(_T_2325_14) : $signed(_GEN_494);
  assign _GEN_496 = 4'hf == _T_1853 ? $signed(_T_2325_15) : $signed(_GEN_495);
  assign _GEN_31 = _GEN_511;
  assign _GEN_497 = 4'h1 == _T_1854 ? $signed(_T_2395_1) : $signed(_T_2395_0);
  assign _GEN_498 = 4'h2 == _T_1854 ? $signed(_T_2395_2) : $signed(_GEN_497);
  assign _GEN_499 = 4'h3 == _T_1854 ? $signed(_T_2395_3) : $signed(_GEN_498);
  assign _GEN_500 = 4'h4 == _T_1854 ? $signed(_T_2395_4) : $signed(_GEN_499);
  assign _GEN_501 = 4'h5 == _T_1854 ? $signed(_T_2395_5) : $signed(_GEN_500);
  assign _GEN_502 = 4'h6 == _T_1854 ? $signed(_T_2395_6) : $signed(_GEN_501);
  assign _GEN_503 = 4'h7 == _T_1854 ? $signed(_T_2395_7) : $signed(_GEN_502);
  assign _GEN_504 = 4'h8 == _T_1854 ? $signed(_T_2395_8) : $signed(_GEN_503);
  assign _GEN_505 = 4'h9 == _T_1854 ? $signed(_T_2395_9) : $signed(_GEN_504);
  assign _GEN_506 = 4'ha == _T_1854 ? $signed(_T_2395_10) : $signed(_GEN_505);
  assign _GEN_507 = 4'hb == _T_1854 ? $signed(_T_2395_11) : $signed(_GEN_506);
  assign _GEN_508 = 4'hc == _T_1854 ? $signed(_T_2395_12) : $signed(_GEN_507);
  assign _GEN_509 = 4'hd == _T_1854 ? $signed(_T_2395_13) : $signed(_GEN_508);
  assign _GEN_510 = 4'he == _T_1854 ? $signed(_T_2395_14) : $signed(_GEN_509);
  assign _GEN_511 = 4'hf == _T_1854 ? $signed(_T_2395_15) : $signed(_GEN_510);
  assign _T_2424 = $signed(_GEN_30) + $signed(_GEN_31);
  assign _T_2425 = _T_2424[5:0];
  assign _T_2426 = $signed(_T_2425);
  assign _T_2427 = $signed(_T_2417) + $signed(_T_2420);
  assign _T_2428 = _T_2427[5:0];
  assign _T_2429 = $signed(_T_2428);
  assign _T_2430 = $signed(_T_2423) + $signed(_T_2426);
  assign _T_2431 = _T_2430[5:0];
  assign _T_2432 = $signed(_T_2431);
  assign _T_2433 = $signed(_T_2429) + $signed(_T_2432);
  assign _T_2434 = _T_2433[5:0];
  assign _T_2435 = $signed(_T_2434);
  assign MulAdd_3_io_a = _T_2438;
  assign MulAdd_3_io_b = Accumulator_3_io_out;
  assign MulAdd_3_io_m = mean_io_output;
  assign MulAdd_3_io_c = _T_2440;
  assign _T_2436 = mem_io_out[31:0];
  assign _T_2437 = _T_2436[31:16];
  assign _T_2438 = $signed(_T_2437);
  assign _T_2439 = _T_2436[15:0];
  assign _T_2440 = $signed(_T_2439);
  assign _T_2441 = MulAdd_3_io_r[31];
  assign signs_3 = ~ _T_2441;
  assign _T_2442 = {signs_2,signs_3};
  assign _T_2443 = {signs_0,signs_1};
  assign _T_2444 = {_T_2443,_T_2442};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_518 = {1{$random}};
  _T_72 = _GEN_518[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_519 = {1{$random}};
  _T_75 = _GEN_519[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_520 = {1{$random}};
  _T_78 = _GEN_520[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_521 = {1{$random}};
  _T_81 = _GEN_521[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_522 = {1{$random}};
  _T_84 = _GEN_522[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_523 = {1{$random}};
  _T_87 = _GEN_523[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_524 = {1{$random}};
  _T_90 = _GEN_524[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_525 = {1{$random}};
  _T_93 = _GEN_525[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_526 = {1{$random}};
  _T_96 = _GEN_526[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_527 = {1{$random}};
  _T_99 = _GEN_527[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_528 = {1{$random}};
  _T_102 = _GEN_528[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_529 = {1{$random}};
  _T_105 = _GEN_529[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_530 = {1{$random}};
  _T_108 = _GEN_530[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_531 = {1{$random}};
  _T_111 = _GEN_531[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_532 = {1{$random}};
  _T_114 = _GEN_532[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_533 = {1{$random}};
  _T_117 = _GEN_533[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_534 = {1{$random}};
  _T_142 = _GEN_534[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_535 = {1{$random}};
  _T_145 = _GEN_535[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_536 = {1{$random}};
  _T_148 = _GEN_536[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_537 = {1{$random}};
  _T_151 = _GEN_537[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_538 = {1{$random}};
  _T_154 = _GEN_538[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_539 = {1{$random}};
  _T_157 = _GEN_539[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_540 = {1{$random}};
  _T_160 = _GEN_540[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_541 = {1{$random}};
  _T_163 = _GEN_541[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_542 = {1{$random}};
  _T_166 = _GEN_542[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_543 = {1{$random}};
  _T_169 = _GEN_543[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_544 = {1{$random}};
  _T_172 = _GEN_544[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_545 = {1{$random}};
  _T_175 = _GEN_545[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_546 = {1{$random}};
  _T_178 = _GEN_546[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_547 = {1{$random}};
  _T_181 = _GEN_547[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_548 = {1{$random}};
  _T_184 = _GEN_548[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_549 = {1{$random}};
  _T_187 = _GEN_549[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_550 = {1{$random}};
  _T_212 = _GEN_550[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_551 = {1{$random}};
  _T_215 = _GEN_551[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_552 = {1{$random}};
  _T_218 = _GEN_552[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_553 = {1{$random}};
  _T_221 = _GEN_553[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_554 = {1{$random}};
  _T_224 = _GEN_554[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_555 = {1{$random}};
  _T_227 = _GEN_555[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_556 = {1{$random}};
  _T_230 = _GEN_556[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_557 = {1{$random}};
  _T_233 = _GEN_557[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_558 = {1{$random}};
  _T_236 = _GEN_558[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_559 = {1{$random}};
  _T_239 = _GEN_559[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_560 = {1{$random}};
  _T_242 = _GEN_560[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_561 = {1{$random}};
  _T_245 = _GEN_561[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_562 = {1{$random}};
  _T_248 = _GEN_562[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_563 = {1{$random}};
  _T_251 = _GEN_563[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_564 = {1{$random}};
  _T_254 = _GEN_564[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_565 = {1{$random}};
  _T_257 = _GEN_565[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_566 = {1{$random}};
  _T_282 = _GEN_566[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_567 = {1{$random}};
  _T_285 = _GEN_567[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_568 = {1{$random}};
  _T_288 = _GEN_568[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_569 = {1{$random}};
  _T_291 = _GEN_569[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_570 = {1{$random}};
  _T_294 = _GEN_570[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_571 = {1{$random}};
  _T_297 = _GEN_571[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_572 = {1{$random}};
  _T_300 = _GEN_572[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_573 = {1{$random}};
  _T_303 = _GEN_573[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_574 = {1{$random}};
  _T_306 = _GEN_574[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_575 = {1{$random}};
  _T_309 = _GEN_575[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_576 = {1{$random}};
  _T_312 = _GEN_576[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_577 = {1{$random}};
  _T_315 = _GEN_577[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_578 = {1{$random}};
  _T_318 = _GEN_578[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_579 = {1{$random}};
  _T_321 = _GEN_579[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_580 = {1{$random}};
  _T_324 = _GEN_580[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_581 = {1{$random}};
  _T_327 = _GEN_581[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_582 = {1{$random}};
  _T_352 = _GEN_582[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_583 = {1{$random}};
  _T_355 = _GEN_583[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_584 = {1{$random}};
  _T_358 = _GEN_584[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_585 = {1{$random}};
  _T_361 = _GEN_585[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_586 = {1{$random}};
  _T_364 = _GEN_586[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_587 = {1{$random}};
  _T_367 = _GEN_587[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_588 = {1{$random}};
  _T_370 = _GEN_588[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_589 = {1{$random}};
  _T_373 = _GEN_589[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_590 = {1{$random}};
  _T_376 = _GEN_590[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_591 = {1{$random}};
  _T_379 = _GEN_591[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_592 = {1{$random}};
  _T_382 = _GEN_592[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_593 = {1{$random}};
  _T_385 = _GEN_593[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_594 = {1{$random}};
  _T_388 = _GEN_594[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_595 = {1{$random}};
  _T_391 = _GEN_595[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_596 = {1{$random}};
  _T_394 = _GEN_596[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_597 = {1{$random}};
  _T_397 = _GEN_597[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_598 = {1{$random}};
  _T_422 = _GEN_598[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_599 = {1{$random}};
  _T_425 = _GEN_599[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_600 = {1{$random}};
  _T_428 = _GEN_600[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_601 = {1{$random}};
  _T_431 = _GEN_601[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_602 = {1{$random}};
  _T_434 = _GEN_602[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_603 = {1{$random}};
  _T_437 = _GEN_603[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_604 = {1{$random}};
  _T_440 = _GEN_604[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_605 = {1{$random}};
  _T_443 = _GEN_605[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_606 = {1{$random}};
  _T_446 = _GEN_606[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_607 = {1{$random}};
  _T_449 = _GEN_607[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_608 = {1{$random}};
  _T_452 = _GEN_608[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_609 = {1{$random}};
  _T_455 = _GEN_609[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_610 = {1{$random}};
  _T_458 = _GEN_610[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_611 = {1{$random}};
  _T_461 = _GEN_611[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_612 = {1{$random}};
  _T_464 = _GEN_612[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_613 = {1{$random}};
  _T_467 = _GEN_613[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_614 = {1{$random}};
  _T_492 = _GEN_614[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_615 = {1{$random}};
  _T_495 = _GEN_615[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_616 = {1{$random}};
  _T_498 = _GEN_616[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_617 = {1{$random}};
  _T_501 = _GEN_617[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_618 = {1{$random}};
  _T_504 = _GEN_618[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_619 = {1{$random}};
  _T_507 = _GEN_619[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_620 = {1{$random}};
  _T_510 = _GEN_620[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_621 = {1{$random}};
  _T_513 = _GEN_621[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_622 = {1{$random}};
  _T_516 = _GEN_622[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_623 = {1{$random}};
  _T_519 = _GEN_623[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_624 = {1{$random}};
  _T_522 = _GEN_624[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_625 = {1{$random}};
  _T_525 = _GEN_625[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_626 = {1{$random}};
  _T_528 = _GEN_626[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_627 = {1{$random}};
  _T_531 = _GEN_627[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_628 = {1{$random}};
  _T_534 = _GEN_628[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_629 = {1{$random}};
  _T_537 = _GEN_629[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_630 = {1{$random}};
  _T_562 = _GEN_630[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_631 = {1{$random}};
  _T_565 = _GEN_631[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_632 = {1{$random}};
  _T_568 = _GEN_632[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_633 = {1{$random}};
  _T_571 = _GEN_633[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_634 = {1{$random}};
  _T_574 = _GEN_634[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_635 = {1{$random}};
  _T_577 = _GEN_635[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_636 = {1{$random}};
  _T_580 = _GEN_636[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_637 = {1{$random}};
  _T_583 = _GEN_637[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_638 = {1{$random}};
  _T_586 = _GEN_638[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_639 = {1{$random}};
  _T_589 = _GEN_639[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_640 = {1{$random}};
  _T_592 = _GEN_640[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_641 = {1{$random}};
  _T_595 = _GEN_641[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_642 = {1{$random}};
  _T_598 = _GEN_642[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_643 = {1{$random}};
  _T_601 = _GEN_643[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_644 = {1{$random}};
  _T_604 = _GEN_644[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_645 = {1{$random}};
  _T_607 = _GEN_645[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_646 = {1{$random}};
  _T_667 = _GEN_646[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_647 = {1{$random}};
  _T_670 = _GEN_647[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_648 = {1{$random}};
  _T_673 = _GEN_648[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_649 = {1{$random}};
  _T_676 = _GEN_649[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_650 = {1{$random}};
  _T_679 = _GEN_650[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_651 = {1{$random}};
  _T_682 = _GEN_651[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_652 = {1{$random}};
  _T_685 = _GEN_652[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_653 = {1{$random}};
  _T_688 = _GEN_653[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_654 = {1{$random}};
  _T_691 = _GEN_654[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_655 = {1{$random}};
  _T_694 = _GEN_655[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_656 = {1{$random}};
  _T_697 = _GEN_656[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_657 = {1{$random}};
  _T_700 = _GEN_657[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_658 = {1{$random}};
  _T_703 = _GEN_658[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_659 = {1{$random}};
  _T_706 = _GEN_659[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_660 = {1{$random}};
  _T_709 = _GEN_660[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_661 = {1{$random}};
  _T_712 = _GEN_661[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_662 = {1{$random}};
  _T_737 = _GEN_662[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_663 = {1{$random}};
  _T_740 = _GEN_663[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_664 = {1{$random}};
  _T_743 = _GEN_664[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_665 = {1{$random}};
  _T_746 = _GEN_665[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_666 = {1{$random}};
  _T_749 = _GEN_666[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_667 = {1{$random}};
  _T_752 = _GEN_667[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_668 = {1{$random}};
  _T_755 = _GEN_668[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_669 = {1{$random}};
  _T_758 = _GEN_669[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_670 = {1{$random}};
  _T_761 = _GEN_670[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_671 = {1{$random}};
  _T_764 = _GEN_671[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_672 = {1{$random}};
  _T_767 = _GEN_672[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_673 = {1{$random}};
  _T_770 = _GEN_673[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_674 = {1{$random}};
  _T_773 = _GEN_674[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_675 = {1{$random}};
  _T_776 = _GEN_675[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_676 = {1{$random}};
  _T_779 = _GEN_676[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_677 = {1{$random}};
  _T_782 = _GEN_677[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_678 = {1{$random}};
  _T_807 = _GEN_678[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_679 = {1{$random}};
  _T_810 = _GEN_679[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_680 = {1{$random}};
  _T_813 = _GEN_680[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_681 = {1{$random}};
  _T_816 = _GEN_681[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_682 = {1{$random}};
  _T_819 = _GEN_682[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_683 = {1{$random}};
  _T_822 = _GEN_683[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_684 = {1{$random}};
  _T_825 = _GEN_684[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_685 = {1{$random}};
  _T_828 = _GEN_685[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_686 = {1{$random}};
  _T_831 = _GEN_686[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_687 = {1{$random}};
  _T_834 = _GEN_687[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_688 = {1{$random}};
  _T_837 = _GEN_688[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_689 = {1{$random}};
  _T_840 = _GEN_689[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_690 = {1{$random}};
  _T_843 = _GEN_690[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_691 = {1{$random}};
  _T_846 = _GEN_691[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_692 = {1{$random}};
  _T_849 = _GEN_692[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_693 = {1{$random}};
  _T_852 = _GEN_693[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_694 = {1{$random}};
  _T_877 = _GEN_694[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_695 = {1{$random}};
  _T_880 = _GEN_695[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_696 = {1{$random}};
  _T_883 = _GEN_696[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_697 = {1{$random}};
  _T_886 = _GEN_697[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_698 = {1{$random}};
  _T_889 = _GEN_698[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_699 = {1{$random}};
  _T_892 = _GEN_699[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_700 = {1{$random}};
  _T_895 = _GEN_700[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_701 = {1{$random}};
  _T_898 = _GEN_701[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_702 = {1{$random}};
  _T_901 = _GEN_702[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_703 = {1{$random}};
  _T_904 = _GEN_703[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_704 = {1{$random}};
  _T_907 = _GEN_704[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_705 = {1{$random}};
  _T_910 = _GEN_705[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_706 = {1{$random}};
  _T_913 = _GEN_706[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_707 = {1{$random}};
  _T_916 = _GEN_707[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_708 = {1{$random}};
  _T_919 = _GEN_708[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_709 = {1{$random}};
  _T_922 = _GEN_709[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_710 = {1{$random}};
  _T_947 = _GEN_710[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_711 = {1{$random}};
  _T_950 = _GEN_711[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_712 = {1{$random}};
  _T_953 = _GEN_712[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_713 = {1{$random}};
  _T_956 = _GEN_713[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_714 = {1{$random}};
  _T_959 = _GEN_714[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_715 = {1{$random}};
  _T_962 = _GEN_715[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_716 = {1{$random}};
  _T_965 = _GEN_716[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_717 = {1{$random}};
  _T_968 = _GEN_717[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_718 = {1{$random}};
  _T_971 = _GEN_718[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_719 = {1{$random}};
  _T_974 = _GEN_719[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_720 = {1{$random}};
  _T_977 = _GEN_720[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_721 = {1{$random}};
  _T_980 = _GEN_721[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_722 = {1{$random}};
  _T_983 = _GEN_722[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_723 = {1{$random}};
  _T_986 = _GEN_723[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_724 = {1{$random}};
  _T_989 = _GEN_724[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_725 = {1{$random}};
  _T_992 = _GEN_725[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_726 = {1{$random}};
  _T_1017 = _GEN_726[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_727 = {1{$random}};
  _T_1020 = _GEN_727[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_728 = {1{$random}};
  _T_1023 = _GEN_728[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_729 = {1{$random}};
  _T_1026 = _GEN_729[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_730 = {1{$random}};
  _T_1029 = _GEN_730[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_731 = {1{$random}};
  _T_1032 = _GEN_731[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_732 = {1{$random}};
  _T_1035 = _GEN_732[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_733 = {1{$random}};
  _T_1038 = _GEN_733[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_734 = {1{$random}};
  _T_1041 = _GEN_734[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_735 = {1{$random}};
  _T_1044 = _GEN_735[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_736 = {1{$random}};
  _T_1047 = _GEN_736[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_737 = {1{$random}};
  _T_1050 = _GEN_737[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_738 = {1{$random}};
  _T_1053 = _GEN_738[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_739 = {1{$random}};
  _T_1056 = _GEN_739[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_740 = {1{$random}};
  _T_1059 = _GEN_740[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_741 = {1{$random}};
  _T_1062 = _GEN_741[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_742 = {1{$random}};
  _T_1087 = _GEN_742[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_743 = {1{$random}};
  _T_1090 = _GEN_743[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_744 = {1{$random}};
  _T_1093 = _GEN_744[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_745 = {1{$random}};
  _T_1096 = _GEN_745[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_746 = {1{$random}};
  _T_1099 = _GEN_746[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_747 = {1{$random}};
  _T_1102 = _GEN_747[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_748 = {1{$random}};
  _T_1105 = _GEN_748[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_749 = {1{$random}};
  _T_1108 = _GEN_749[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_750 = {1{$random}};
  _T_1111 = _GEN_750[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_751 = {1{$random}};
  _T_1114 = _GEN_751[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_752 = {1{$random}};
  _T_1117 = _GEN_752[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_753 = {1{$random}};
  _T_1120 = _GEN_753[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_754 = {1{$random}};
  _T_1123 = _GEN_754[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_755 = {1{$random}};
  _T_1126 = _GEN_755[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_756 = {1{$random}};
  _T_1129 = _GEN_756[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_757 = {1{$random}};
  _T_1132 = _GEN_757[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_758 = {1{$random}};
  _T_1157 = _GEN_758[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_759 = {1{$random}};
  _T_1160 = _GEN_759[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_760 = {1{$random}};
  _T_1163 = _GEN_760[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_761 = {1{$random}};
  _T_1166 = _GEN_761[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_762 = {1{$random}};
  _T_1169 = _GEN_762[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_763 = {1{$random}};
  _T_1172 = _GEN_763[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_764 = {1{$random}};
  _T_1175 = _GEN_764[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_765 = {1{$random}};
  _T_1178 = _GEN_765[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_766 = {1{$random}};
  _T_1181 = _GEN_766[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_767 = {1{$random}};
  _T_1184 = _GEN_767[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_768 = {1{$random}};
  _T_1187 = _GEN_768[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_769 = {1{$random}};
  _T_1190 = _GEN_769[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_770 = {1{$random}};
  _T_1193 = _GEN_770[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_771 = {1{$random}};
  _T_1196 = _GEN_771[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_772 = {1{$random}};
  _T_1199 = _GEN_772[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_773 = {1{$random}};
  _T_1202 = _GEN_773[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_774 = {1{$random}};
  _T_1262 = _GEN_774[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_775 = {1{$random}};
  _T_1265 = _GEN_775[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_776 = {1{$random}};
  _T_1268 = _GEN_776[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_777 = {1{$random}};
  _T_1271 = _GEN_777[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_778 = {1{$random}};
  _T_1274 = _GEN_778[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_779 = {1{$random}};
  _T_1277 = _GEN_779[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_780 = {1{$random}};
  _T_1280 = _GEN_780[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_781 = {1{$random}};
  _T_1283 = _GEN_781[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_782 = {1{$random}};
  _T_1286 = _GEN_782[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_783 = {1{$random}};
  _T_1289 = _GEN_783[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_784 = {1{$random}};
  _T_1292 = _GEN_784[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_785 = {1{$random}};
  _T_1295 = _GEN_785[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_786 = {1{$random}};
  _T_1298 = _GEN_786[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_787 = {1{$random}};
  _T_1301 = _GEN_787[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_788 = {1{$random}};
  _T_1304 = _GEN_788[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_789 = {1{$random}};
  _T_1307 = _GEN_789[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_790 = {1{$random}};
  _T_1332 = _GEN_790[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_791 = {1{$random}};
  _T_1335 = _GEN_791[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_792 = {1{$random}};
  _T_1338 = _GEN_792[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_793 = {1{$random}};
  _T_1341 = _GEN_793[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_794 = {1{$random}};
  _T_1344 = _GEN_794[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_795 = {1{$random}};
  _T_1347 = _GEN_795[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_796 = {1{$random}};
  _T_1350 = _GEN_796[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_797 = {1{$random}};
  _T_1353 = _GEN_797[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_798 = {1{$random}};
  _T_1356 = _GEN_798[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_799 = {1{$random}};
  _T_1359 = _GEN_799[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_800 = {1{$random}};
  _T_1362 = _GEN_800[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_801 = {1{$random}};
  _T_1365 = _GEN_801[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_802 = {1{$random}};
  _T_1368 = _GEN_802[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_803 = {1{$random}};
  _T_1371 = _GEN_803[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_804 = {1{$random}};
  _T_1374 = _GEN_804[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_805 = {1{$random}};
  _T_1377 = _GEN_805[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_806 = {1{$random}};
  _T_1402 = _GEN_806[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_807 = {1{$random}};
  _T_1405 = _GEN_807[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_808 = {1{$random}};
  _T_1408 = _GEN_808[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_809 = {1{$random}};
  _T_1411 = _GEN_809[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_810 = {1{$random}};
  _T_1414 = _GEN_810[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_811 = {1{$random}};
  _T_1417 = _GEN_811[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_812 = {1{$random}};
  _T_1420 = _GEN_812[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_813 = {1{$random}};
  _T_1423 = _GEN_813[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_814 = {1{$random}};
  _T_1426 = _GEN_814[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_815 = {1{$random}};
  _T_1429 = _GEN_815[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_816 = {1{$random}};
  _T_1432 = _GEN_816[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_817 = {1{$random}};
  _T_1435 = _GEN_817[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_818 = {1{$random}};
  _T_1438 = _GEN_818[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_819 = {1{$random}};
  _T_1441 = _GEN_819[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_820 = {1{$random}};
  _T_1444 = _GEN_820[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_821 = {1{$random}};
  _T_1447 = _GEN_821[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_822 = {1{$random}};
  _T_1472 = _GEN_822[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_823 = {1{$random}};
  _T_1475 = _GEN_823[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_824 = {1{$random}};
  _T_1478 = _GEN_824[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_825 = {1{$random}};
  _T_1481 = _GEN_825[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_826 = {1{$random}};
  _T_1484 = _GEN_826[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_827 = {1{$random}};
  _T_1487 = _GEN_827[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_828 = {1{$random}};
  _T_1490 = _GEN_828[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_829 = {1{$random}};
  _T_1493 = _GEN_829[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_830 = {1{$random}};
  _T_1496 = _GEN_830[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_831 = {1{$random}};
  _T_1499 = _GEN_831[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_832 = {1{$random}};
  _T_1502 = _GEN_832[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_833 = {1{$random}};
  _T_1505 = _GEN_833[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_834 = {1{$random}};
  _T_1508 = _GEN_834[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_835 = {1{$random}};
  _T_1511 = _GEN_835[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_836 = {1{$random}};
  _T_1514 = _GEN_836[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_837 = {1{$random}};
  _T_1517 = _GEN_837[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_838 = {1{$random}};
  _T_1542 = _GEN_838[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_839 = {1{$random}};
  _T_1545 = _GEN_839[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_840 = {1{$random}};
  _T_1548 = _GEN_840[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_841 = {1{$random}};
  _T_1551 = _GEN_841[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_842 = {1{$random}};
  _T_1554 = _GEN_842[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_843 = {1{$random}};
  _T_1557 = _GEN_843[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_844 = {1{$random}};
  _T_1560 = _GEN_844[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_845 = {1{$random}};
  _T_1563 = _GEN_845[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_846 = {1{$random}};
  _T_1566 = _GEN_846[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_847 = {1{$random}};
  _T_1569 = _GEN_847[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_848 = {1{$random}};
  _T_1572 = _GEN_848[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_849 = {1{$random}};
  _T_1575 = _GEN_849[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_850 = {1{$random}};
  _T_1578 = _GEN_850[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_851 = {1{$random}};
  _T_1581 = _GEN_851[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_852 = {1{$random}};
  _T_1584 = _GEN_852[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_853 = {1{$random}};
  _T_1587 = _GEN_853[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_854 = {1{$random}};
  _T_1612 = _GEN_854[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_855 = {1{$random}};
  _T_1615 = _GEN_855[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_856 = {1{$random}};
  _T_1618 = _GEN_856[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_857 = {1{$random}};
  _T_1621 = _GEN_857[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_858 = {1{$random}};
  _T_1624 = _GEN_858[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_859 = {1{$random}};
  _T_1627 = _GEN_859[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_860 = {1{$random}};
  _T_1630 = _GEN_860[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_861 = {1{$random}};
  _T_1633 = _GEN_861[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_862 = {1{$random}};
  _T_1636 = _GEN_862[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_863 = {1{$random}};
  _T_1639 = _GEN_863[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_864 = {1{$random}};
  _T_1642 = _GEN_864[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_865 = {1{$random}};
  _T_1645 = _GEN_865[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_866 = {1{$random}};
  _T_1648 = _GEN_866[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_867 = {1{$random}};
  _T_1651 = _GEN_867[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_868 = {1{$random}};
  _T_1654 = _GEN_868[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_869 = {1{$random}};
  _T_1657 = _GEN_869[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_870 = {1{$random}};
  _T_1682 = _GEN_870[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_871 = {1{$random}};
  _T_1685 = _GEN_871[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_872 = {1{$random}};
  _T_1688 = _GEN_872[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_873 = {1{$random}};
  _T_1691 = _GEN_873[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_874 = {1{$random}};
  _T_1694 = _GEN_874[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_875 = {1{$random}};
  _T_1697 = _GEN_875[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_876 = {1{$random}};
  _T_1700 = _GEN_876[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_877 = {1{$random}};
  _T_1703 = _GEN_877[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_878 = {1{$random}};
  _T_1706 = _GEN_878[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_879 = {1{$random}};
  _T_1709 = _GEN_879[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_880 = {1{$random}};
  _T_1712 = _GEN_880[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_881 = {1{$random}};
  _T_1715 = _GEN_881[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_882 = {1{$random}};
  _T_1718 = _GEN_882[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_883 = {1{$random}};
  _T_1721 = _GEN_883[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_884 = {1{$random}};
  _T_1724 = _GEN_884[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_885 = {1{$random}};
  _T_1727 = _GEN_885[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_886 = {1{$random}};
  _T_1752 = _GEN_886[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_887 = {1{$random}};
  _T_1755 = _GEN_887[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_888 = {1{$random}};
  _T_1758 = _GEN_888[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_889 = {1{$random}};
  _T_1761 = _GEN_889[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_890 = {1{$random}};
  _T_1764 = _GEN_890[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_891 = {1{$random}};
  _T_1767 = _GEN_891[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_892 = {1{$random}};
  _T_1770 = _GEN_892[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_893 = {1{$random}};
  _T_1773 = _GEN_893[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_894 = {1{$random}};
  _T_1776 = _GEN_894[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_895 = {1{$random}};
  _T_1779 = _GEN_895[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_896 = {1{$random}};
  _T_1782 = _GEN_896[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_897 = {1{$random}};
  _T_1785 = _GEN_897[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_898 = {1{$random}};
  _T_1788 = _GEN_898[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_899 = {1{$random}};
  _T_1791 = _GEN_899[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_900 = {1{$random}};
  _T_1794 = _GEN_900[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_901 = {1{$random}};
  _T_1797 = _GEN_901[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_902 = {1{$random}};
  _T_1857 = _GEN_902[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_903 = {1{$random}};
  _T_1860 = _GEN_903[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_904 = {1{$random}};
  _T_1863 = _GEN_904[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_905 = {1{$random}};
  _T_1866 = _GEN_905[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_906 = {1{$random}};
  _T_1869 = _GEN_906[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_907 = {1{$random}};
  _T_1872 = _GEN_907[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_908 = {1{$random}};
  _T_1875 = _GEN_908[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_909 = {1{$random}};
  _T_1878 = _GEN_909[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_910 = {1{$random}};
  _T_1881 = _GEN_910[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_911 = {1{$random}};
  _T_1884 = _GEN_911[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_912 = {1{$random}};
  _T_1887 = _GEN_912[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_913 = {1{$random}};
  _T_1890 = _GEN_913[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_914 = {1{$random}};
  _T_1893 = _GEN_914[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_915 = {1{$random}};
  _T_1896 = _GEN_915[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_916 = {1{$random}};
  _T_1899 = _GEN_916[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_917 = {1{$random}};
  _T_1902 = _GEN_917[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_918 = {1{$random}};
  _T_1927 = _GEN_918[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_919 = {1{$random}};
  _T_1930 = _GEN_919[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_920 = {1{$random}};
  _T_1933 = _GEN_920[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_921 = {1{$random}};
  _T_1936 = _GEN_921[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_922 = {1{$random}};
  _T_1939 = _GEN_922[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_923 = {1{$random}};
  _T_1942 = _GEN_923[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_924 = {1{$random}};
  _T_1945 = _GEN_924[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_925 = {1{$random}};
  _T_1948 = _GEN_925[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_926 = {1{$random}};
  _T_1951 = _GEN_926[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_927 = {1{$random}};
  _T_1954 = _GEN_927[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_928 = {1{$random}};
  _T_1957 = _GEN_928[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_929 = {1{$random}};
  _T_1960 = _GEN_929[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_930 = {1{$random}};
  _T_1963 = _GEN_930[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_931 = {1{$random}};
  _T_1966 = _GEN_931[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_932 = {1{$random}};
  _T_1969 = _GEN_932[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_933 = {1{$random}};
  _T_1972 = _GEN_933[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_934 = {1{$random}};
  _T_1997 = _GEN_934[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_935 = {1{$random}};
  _T_2000 = _GEN_935[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_936 = {1{$random}};
  _T_2003 = _GEN_936[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_937 = {1{$random}};
  _T_2006 = _GEN_937[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_938 = {1{$random}};
  _T_2009 = _GEN_938[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_939 = {1{$random}};
  _T_2012 = _GEN_939[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_940 = {1{$random}};
  _T_2015 = _GEN_940[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_941 = {1{$random}};
  _T_2018 = _GEN_941[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_942 = {1{$random}};
  _T_2021 = _GEN_942[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_943 = {1{$random}};
  _T_2024 = _GEN_943[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_944 = {1{$random}};
  _T_2027 = _GEN_944[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_945 = {1{$random}};
  _T_2030 = _GEN_945[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_946 = {1{$random}};
  _T_2033 = _GEN_946[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_947 = {1{$random}};
  _T_2036 = _GEN_947[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_948 = {1{$random}};
  _T_2039 = _GEN_948[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_949 = {1{$random}};
  _T_2042 = _GEN_949[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_950 = {1{$random}};
  _T_2067 = _GEN_950[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_951 = {1{$random}};
  _T_2070 = _GEN_951[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_952 = {1{$random}};
  _T_2073 = _GEN_952[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_953 = {1{$random}};
  _T_2076 = _GEN_953[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_954 = {1{$random}};
  _T_2079 = _GEN_954[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_955 = {1{$random}};
  _T_2082 = _GEN_955[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_956 = {1{$random}};
  _T_2085 = _GEN_956[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_957 = {1{$random}};
  _T_2088 = _GEN_957[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_958 = {1{$random}};
  _T_2091 = _GEN_958[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_959 = {1{$random}};
  _T_2094 = _GEN_959[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_960 = {1{$random}};
  _T_2097 = _GEN_960[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_961 = {1{$random}};
  _T_2100 = _GEN_961[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_962 = {1{$random}};
  _T_2103 = _GEN_962[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_963 = {1{$random}};
  _T_2106 = _GEN_963[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_964 = {1{$random}};
  _T_2109 = _GEN_964[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_965 = {1{$random}};
  _T_2112 = _GEN_965[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_966 = {1{$random}};
  _T_2137 = _GEN_966[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_967 = {1{$random}};
  _T_2140 = _GEN_967[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_968 = {1{$random}};
  _T_2143 = _GEN_968[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_969 = {1{$random}};
  _T_2146 = _GEN_969[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_970 = {1{$random}};
  _T_2149 = _GEN_970[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_971 = {1{$random}};
  _T_2152 = _GEN_971[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_972 = {1{$random}};
  _T_2155 = _GEN_972[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_973 = {1{$random}};
  _T_2158 = _GEN_973[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_974 = {1{$random}};
  _T_2161 = _GEN_974[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_975 = {1{$random}};
  _T_2164 = _GEN_975[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_976 = {1{$random}};
  _T_2167 = _GEN_976[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_977 = {1{$random}};
  _T_2170 = _GEN_977[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_978 = {1{$random}};
  _T_2173 = _GEN_978[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_979 = {1{$random}};
  _T_2176 = _GEN_979[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_980 = {1{$random}};
  _T_2179 = _GEN_980[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_981 = {1{$random}};
  _T_2182 = _GEN_981[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_982 = {1{$random}};
  _T_2207 = _GEN_982[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_983 = {1{$random}};
  _T_2210 = _GEN_983[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_984 = {1{$random}};
  _T_2213 = _GEN_984[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_985 = {1{$random}};
  _T_2216 = _GEN_985[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_986 = {1{$random}};
  _T_2219 = _GEN_986[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_987 = {1{$random}};
  _T_2222 = _GEN_987[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_988 = {1{$random}};
  _T_2225 = _GEN_988[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_989 = {1{$random}};
  _T_2228 = _GEN_989[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_990 = {1{$random}};
  _T_2231 = _GEN_990[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_991 = {1{$random}};
  _T_2234 = _GEN_991[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_992 = {1{$random}};
  _T_2237 = _GEN_992[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_993 = {1{$random}};
  _T_2240 = _GEN_993[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_994 = {1{$random}};
  _T_2243 = _GEN_994[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_995 = {1{$random}};
  _T_2246 = _GEN_995[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_996 = {1{$random}};
  _T_2249 = _GEN_996[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_997 = {1{$random}};
  _T_2252 = _GEN_997[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_998 = {1{$random}};
  _T_2277 = _GEN_998[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_999 = {1{$random}};
  _T_2280 = _GEN_999[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1000 = {1{$random}};
  _T_2283 = _GEN_1000[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1001 = {1{$random}};
  _T_2286 = _GEN_1001[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1002 = {1{$random}};
  _T_2289 = _GEN_1002[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1003 = {1{$random}};
  _T_2292 = _GEN_1003[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1004 = {1{$random}};
  _T_2295 = _GEN_1004[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1005 = {1{$random}};
  _T_2298 = _GEN_1005[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1006 = {1{$random}};
  _T_2301 = _GEN_1006[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1007 = {1{$random}};
  _T_2304 = _GEN_1007[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1008 = {1{$random}};
  _T_2307 = _GEN_1008[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1009 = {1{$random}};
  _T_2310 = _GEN_1009[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1010 = {1{$random}};
  _T_2313 = _GEN_1010[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1011 = {1{$random}};
  _T_2316 = _GEN_1011[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1012 = {1{$random}};
  _T_2319 = _GEN_1012[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1013 = {1{$random}};
  _T_2322 = _GEN_1013[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1014 = {1{$random}};
  _T_2347 = _GEN_1014[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1015 = {1{$random}};
  _T_2350 = _GEN_1015[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1016 = {1{$random}};
  _T_2353 = _GEN_1016[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1017 = {1{$random}};
  _T_2356 = _GEN_1017[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1018 = {1{$random}};
  _T_2359 = _GEN_1018[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1019 = {1{$random}};
  _T_2362 = _GEN_1019[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1020 = {1{$random}};
  _T_2365 = _GEN_1020[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1021 = {1{$random}};
  _T_2368 = _GEN_1021[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1022 = {1{$random}};
  _T_2371 = _GEN_1022[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1023 = {1{$random}};
  _T_2374 = _GEN_1023[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1024 = {1{$random}};
  _T_2377 = _GEN_1024[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1025 = {1{$random}};
  _T_2380 = _GEN_1025[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1026 = {1{$random}};
  _T_2383 = _GEN_1026[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1027 = {1{$random}};
  _T_2386 = _GEN_1027[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1028 = {1{$random}};
  _T_2389 = _GEN_1028[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1029 = {1{$random}};
  _T_2392 = _GEN_1029[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1030 = {1{$random}};
  _GEN_512 = _GEN_1030[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1031 = {1{$random}};
  _GEN_513 = _GEN_1031[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1032 = {1{$random}};
  _GEN_514 = _GEN_1032[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1033 = {1{$random}};
  _GEN_515 = _GEN_1033[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1034 = {1{$random}};
  _GEN_516 = _GEN_1034[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1035 = {1{$random}};
  _GEN_517 = _GEN_1035[15:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (reset) begin
      _T_72 <= -6'sh4;
    end
    if (reset) begin
      _T_75 <= -6'sh2;
    end
    if (reset) begin
      _T_78 <= -6'sh2;
    end
    if (reset) begin
      _T_81 <= 6'sh0;
    end
    if (reset) begin
      _T_84 <= -6'sh2;
    end
    if (reset) begin
      _T_87 <= 6'sh0;
    end
    if (reset) begin
      _T_90 <= 6'sh0;
    end
    if (reset) begin
      _T_93 <= 6'sh2;
    end
    if (reset) begin
      _T_96 <= -6'sh2;
    end
    if (reset) begin
      _T_99 <= 6'sh0;
    end
    if (reset) begin
      _T_102 <= 6'sh0;
    end
    if (reset) begin
      _T_105 <= 6'sh2;
    end
    if (reset) begin
      _T_108 <= 6'sh0;
    end
    if (reset) begin
      _T_111 <= 6'sh2;
    end
    if (reset) begin
      _T_114 <= 6'sh2;
    end
    if (reset) begin
      _T_117 <= 6'sh4;
    end
    if (reset) begin
      _T_142 <= -6'sh4;
    end
    if (reset) begin
      _T_145 <= -6'sh2;
    end
    if (reset) begin
      _T_148 <= -6'sh2;
    end
    if (reset) begin
      _T_151 <= 6'sh0;
    end
    if (reset) begin
      _T_154 <= -6'sh2;
    end
    if (reset) begin
      _T_157 <= 6'sh0;
    end
    if (reset) begin
      _T_160 <= 6'sh0;
    end
    if (reset) begin
      _T_163 <= 6'sh2;
    end
    if (reset) begin
      _T_166 <= -6'sh2;
    end
    if (reset) begin
      _T_169 <= 6'sh0;
    end
    if (reset) begin
      _T_172 <= 6'sh0;
    end
    if (reset) begin
      _T_175 <= 6'sh2;
    end
    if (reset) begin
      _T_178 <= 6'sh0;
    end
    if (reset) begin
      _T_181 <= 6'sh2;
    end
    if (reset) begin
      _T_184 <= 6'sh2;
    end
    if (reset) begin
      _T_187 <= 6'sh4;
    end
    if (reset) begin
      _T_212 <= -6'sh4;
    end
    if (reset) begin
      _T_215 <= -6'sh2;
    end
    if (reset) begin
      _T_218 <= -6'sh2;
    end
    if (reset) begin
      _T_221 <= 6'sh0;
    end
    if (reset) begin
      _T_224 <= -6'sh2;
    end
    if (reset) begin
      _T_227 <= 6'sh0;
    end
    if (reset) begin
      _T_230 <= 6'sh0;
    end
    if (reset) begin
      _T_233 <= 6'sh2;
    end
    if (reset) begin
      _T_236 <= -6'sh2;
    end
    if (reset) begin
      _T_239 <= 6'sh0;
    end
    if (reset) begin
      _T_242 <= 6'sh0;
    end
    if (reset) begin
      _T_245 <= 6'sh2;
    end
    if (reset) begin
      _T_248 <= 6'sh0;
    end
    if (reset) begin
      _T_251 <= 6'sh2;
    end
    if (reset) begin
      _T_254 <= 6'sh2;
    end
    if (reset) begin
      _T_257 <= 6'sh4;
    end
    if (reset) begin
      _T_282 <= -6'sh4;
    end
    if (reset) begin
      _T_285 <= -6'sh2;
    end
    if (reset) begin
      _T_288 <= -6'sh2;
    end
    if (reset) begin
      _T_291 <= 6'sh0;
    end
    if (reset) begin
      _T_294 <= -6'sh2;
    end
    if (reset) begin
      _T_297 <= 6'sh0;
    end
    if (reset) begin
      _T_300 <= 6'sh0;
    end
    if (reset) begin
      _T_303 <= 6'sh2;
    end
    if (reset) begin
      _T_306 <= -6'sh2;
    end
    if (reset) begin
      _T_309 <= 6'sh0;
    end
    if (reset) begin
      _T_312 <= 6'sh0;
    end
    if (reset) begin
      _T_315 <= 6'sh2;
    end
    if (reset) begin
      _T_318 <= 6'sh0;
    end
    if (reset) begin
      _T_321 <= 6'sh2;
    end
    if (reset) begin
      _T_324 <= 6'sh2;
    end
    if (reset) begin
      _T_327 <= 6'sh4;
    end
    if (reset) begin
      _T_352 <= -6'sh4;
    end
    if (reset) begin
      _T_355 <= -6'sh2;
    end
    if (reset) begin
      _T_358 <= -6'sh2;
    end
    if (reset) begin
      _T_361 <= 6'sh0;
    end
    if (reset) begin
      _T_364 <= -6'sh2;
    end
    if (reset) begin
      _T_367 <= 6'sh0;
    end
    if (reset) begin
      _T_370 <= 6'sh0;
    end
    if (reset) begin
      _T_373 <= 6'sh2;
    end
    if (reset) begin
      _T_376 <= -6'sh2;
    end
    if (reset) begin
      _T_379 <= 6'sh0;
    end
    if (reset) begin
      _T_382 <= 6'sh0;
    end
    if (reset) begin
      _T_385 <= 6'sh2;
    end
    if (reset) begin
      _T_388 <= 6'sh0;
    end
    if (reset) begin
      _T_391 <= 6'sh2;
    end
    if (reset) begin
      _T_394 <= 6'sh2;
    end
    if (reset) begin
      _T_397 <= 6'sh4;
    end
    if (reset) begin
      _T_422 <= -6'sh4;
    end
    if (reset) begin
      _T_425 <= -6'sh2;
    end
    if (reset) begin
      _T_428 <= -6'sh2;
    end
    if (reset) begin
      _T_431 <= 6'sh0;
    end
    if (reset) begin
      _T_434 <= -6'sh2;
    end
    if (reset) begin
      _T_437 <= 6'sh0;
    end
    if (reset) begin
      _T_440 <= 6'sh0;
    end
    if (reset) begin
      _T_443 <= 6'sh2;
    end
    if (reset) begin
      _T_446 <= -6'sh2;
    end
    if (reset) begin
      _T_449 <= 6'sh0;
    end
    if (reset) begin
      _T_452 <= 6'sh0;
    end
    if (reset) begin
      _T_455 <= 6'sh2;
    end
    if (reset) begin
      _T_458 <= 6'sh0;
    end
    if (reset) begin
      _T_461 <= 6'sh2;
    end
    if (reset) begin
      _T_464 <= 6'sh2;
    end
    if (reset) begin
      _T_467 <= 6'sh4;
    end
    if (reset) begin
      _T_492 <= -6'sh4;
    end
    if (reset) begin
      _T_495 <= -6'sh2;
    end
    if (reset) begin
      _T_498 <= -6'sh2;
    end
    if (reset) begin
      _T_501 <= 6'sh0;
    end
    if (reset) begin
      _T_504 <= -6'sh2;
    end
    if (reset) begin
      _T_507 <= 6'sh0;
    end
    if (reset) begin
      _T_510 <= 6'sh0;
    end
    if (reset) begin
      _T_513 <= 6'sh2;
    end
    if (reset) begin
      _T_516 <= -6'sh2;
    end
    if (reset) begin
      _T_519 <= 6'sh0;
    end
    if (reset) begin
      _T_522 <= 6'sh0;
    end
    if (reset) begin
      _T_525 <= 6'sh2;
    end
    if (reset) begin
      _T_528 <= 6'sh0;
    end
    if (reset) begin
      _T_531 <= 6'sh2;
    end
    if (reset) begin
      _T_534 <= 6'sh2;
    end
    if (reset) begin
      _T_537 <= 6'sh4;
    end
    if (reset) begin
      _T_562 <= -6'sh4;
    end
    if (reset) begin
      _T_565 <= -6'sh2;
    end
    if (reset) begin
      _T_568 <= -6'sh2;
    end
    if (reset) begin
      _T_571 <= 6'sh0;
    end
    if (reset) begin
      _T_574 <= -6'sh2;
    end
    if (reset) begin
      _T_577 <= 6'sh0;
    end
    if (reset) begin
      _T_580 <= 6'sh0;
    end
    if (reset) begin
      _T_583 <= 6'sh2;
    end
    if (reset) begin
      _T_586 <= -6'sh2;
    end
    if (reset) begin
      _T_589 <= 6'sh0;
    end
    if (reset) begin
      _T_592 <= 6'sh0;
    end
    if (reset) begin
      _T_595 <= 6'sh2;
    end
    if (reset) begin
      _T_598 <= 6'sh0;
    end
    if (reset) begin
      _T_601 <= 6'sh2;
    end
    if (reset) begin
      _T_604 <= 6'sh2;
    end
    if (reset) begin
      _T_607 <= 6'sh4;
    end
    if (reset) begin
      _T_667 <= -6'sh4;
    end
    if (reset) begin
      _T_670 <= -6'sh2;
    end
    if (reset) begin
      _T_673 <= -6'sh2;
    end
    if (reset) begin
      _T_676 <= 6'sh0;
    end
    if (reset) begin
      _T_679 <= -6'sh2;
    end
    if (reset) begin
      _T_682 <= 6'sh0;
    end
    if (reset) begin
      _T_685 <= 6'sh0;
    end
    if (reset) begin
      _T_688 <= 6'sh2;
    end
    if (reset) begin
      _T_691 <= -6'sh2;
    end
    if (reset) begin
      _T_694 <= 6'sh0;
    end
    if (reset) begin
      _T_697 <= 6'sh0;
    end
    if (reset) begin
      _T_700 <= 6'sh2;
    end
    if (reset) begin
      _T_703 <= 6'sh0;
    end
    if (reset) begin
      _T_706 <= 6'sh2;
    end
    if (reset) begin
      _T_709 <= 6'sh2;
    end
    if (reset) begin
      _T_712 <= 6'sh4;
    end
    if (reset) begin
      _T_737 <= -6'sh4;
    end
    if (reset) begin
      _T_740 <= -6'sh2;
    end
    if (reset) begin
      _T_743 <= -6'sh2;
    end
    if (reset) begin
      _T_746 <= 6'sh0;
    end
    if (reset) begin
      _T_749 <= -6'sh2;
    end
    if (reset) begin
      _T_752 <= 6'sh0;
    end
    if (reset) begin
      _T_755 <= 6'sh0;
    end
    if (reset) begin
      _T_758 <= 6'sh2;
    end
    if (reset) begin
      _T_761 <= -6'sh2;
    end
    if (reset) begin
      _T_764 <= 6'sh0;
    end
    if (reset) begin
      _T_767 <= 6'sh0;
    end
    if (reset) begin
      _T_770 <= 6'sh2;
    end
    if (reset) begin
      _T_773 <= 6'sh0;
    end
    if (reset) begin
      _T_776 <= 6'sh2;
    end
    if (reset) begin
      _T_779 <= 6'sh2;
    end
    if (reset) begin
      _T_782 <= 6'sh4;
    end
    if (reset) begin
      _T_807 <= -6'sh4;
    end
    if (reset) begin
      _T_810 <= -6'sh2;
    end
    if (reset) begin
      _T_813 <= -6'sh2;
    end
    if (reset) begin
      _T_816 <= 6'sh0;
    end
    if (reset) begin
      _T_819 <= -6'sh2;
    end
    if (reset) begin
      _T_822 <= 6'sh0;
    end
    if (reset) begin
      _T_825 <= 6'sh0;
    end
    if (reset) begin
      _T_828 <= 6'sh2;
    end
    if (reset) begin
      _T_831 <= -6'sh2;
    end
    if (reset) begin
      _T_834 <= 6'sh0;
    end
    if (reset) begin
      _T_837 <= 6'sh0;
    end
    if (reset) begin
      _T_840 <= 6'sh2;
    end
    if (reset) begin
      _T_843 <= 6'sh0;
    end
    if (reset) begin
      _T_846 <= 6'sh2;
    end
    if (reset) begin
      _T_849 <= 6'sh2;
    end
    if (reset) begin
      _T_852 <= 6'sh4;
    end
    if (reset) begin
      _T_877 <= -6'sh4;
    end
    if (reset) begin
      _T_880 <= -6'sh2;
    end
    if (reset) begin
      _T_883 <= -6'sh2;
    end
    if (reset) begin
      _T_886 <= 6'sh0;
    end
    if (reset) begin
      _T_889 <= -6'sh2;
    end
    if (reset) begin
      _T_892 <= 6'sh0;
    end
    if (reset) begin
      _T_895 <= 6'sh0;
    end
    if (reset) begin
      _T_898 <= 6'sh2;
    end
    if (reset) begin
      _T_901 <= -6'sh2;
    end
    if (reset) begin
      _T_904 <= 6'sh0;
    end
    if (reset) begin
      _T_907 <= 6'sh0;
    end
    if (reset) begin
      _T_910 <= 6'sh2;
    end
    if (reset) begin
      _T_913 <= 6'sh0;
    end
    if (reset) begin
      _T_916 <= 6'sh2;
    end
    if (reset) begin
      _T_919 <= 6'sh2;
    end
    if (reset) begin
      _T_922 <= 6'sh4;
    end
    if (reset) begin
      _T_947 <= -6'sh4;
    end
    if (reset) begin
      _T_950 <= -6'sh2;
    end
    if (reset) begin
      _T_953 <= -6'sh2;
    end
    if (reset) begin
      _T_956 <= 6'sh0;
    end
    if (reset) begin
      _T_959 <= -6'sh2;
    end
    if (reset) begin
      _T_962 <= 6'sh0;
    end
    if (reset) begin
      _T_965 <= 6'sh0;
    end
    if (reset) begin
      _T_968 <= 6'sh2;
    end
    if (reset) begin
      _T_971 <= -6'sh2;
    end
    if (reset) begin
      _T_974 <= 6'sh0;
    end
    if (reset) begin
      _T_977 <= 6'sh0;
    end
    if (reset) begin
      _T_980 <= 6'sh2;
    end
    if (reset) begin
      _T_983 <= 6'sh0;
    end
    if (reset) begin
      _T_986 <= 6'sh2;
    end
    if (reset) begin
      _T_989 <= 6'sh2;
    end
    if (reset) begin
      _T_992 <= 6'sh4;
    end
    if (reset) begin
      _T_1017 <= -6'sh4;
    end
    if (reset) begin
      _T_1020 <= -6'sh2;
    end
    if (reset) begin
      _T_1023 <= -6'sh2;
    end
    if (reset) begin
      _T_1026 <= 6'sh0;
    end
    if (reset) begin
      _T_1029 <= -6'sh2;
    end
    if (reset) begin
      _T_1032 <= 6'sh0;
    end
    if (reset) begin
      _T_1035 <= 6'sh0;
    end
    if (reset) begin
      _T_1038 <= 6'sh2;
    end
    if (reset) begin
      _T_1041 <= -6'sh2;
    end
    if (reset) begin
      _T_1044 <= 6'sh0;
    end
    if (reset) begin
      _T_1047 <= 6'sh0;
    end
    if (reset) begin
      _T_1050 <= 6'sh2;
    end
    if (reset) begin
      _T_1053 <= 6'sh0;
    end
    if (reset) begin
      _T_1056 <= 6'sh2;
    end
    if (reset) begin
      _T_1059 <= 6'sh2;
    end
    if (reset) begin
      _T_1062 <= 6'sh4;
    end
    if (reset) begin
      _T_1087 <= -6'sh4;
    end
    if (reset) begin
      _T_1090 <= -6'sh2;
    end
    if (reset) begin
      _T_1093 <= -6'sh2;
    end
    if (reset) begin
      _T_1096 <= 6'sh0;
    end
    if (reset) begin
      _T_1099 <= -6'sh2;
    end
    if (reset) begin
      _T_1102 <= 6'sh0;
    end
    if (reset) begin
      _T_1105 <= 6'sh0;
    end
    if (reset) begin
      _T_1108 <= 6'sh2;
    end
    if (reset) begin
      _T_1111 <= -6'sh2;
    end
    if (reset) begin
      _T_1114 <= 6'sh0;
    end
    if (reset) begin
      _T_1117 <= 6'sh0;
    end
    if (reset) begin
      _T_1120 <= 6'sh2;
    end
    if (reset) begin
      _T_1123 <= 6'sh0;
    end
    if (reset) begin
      _T_1126 <= 6'sh2;
    end
    if (reset) begin
      _T_1129 <= 6'sh2;
    end
    if (reset) begin
      _T_1132 <= 6'sh4;
    end
    if (reset) begin
      _T_1157 <= -6'sh4;
    end
    if (reset) begin
      _T_1160 <= -6'sh2;
    end
    if (reset) begin
      _T_1163 <= -6'sh2;
    end
    if (reset) begin
      _T_1166 <= 6'sh0;
    end
    if (reset) begin
      _T_1169 <= -6'sh2;
    end
    if (reset) begin
      _T_1172 <= 6'sh0;
    end
    if (reset) begin
      _T_1175 <= 6'sh0;
    end
    if (reset) begin
      _T_1178 <= 6'sh2;
    end
    if (reset) begin
      _T_1181 <= -6'sh2;
    end
    if (reset) begin
      _T_1184 <= 6'sh0;
    end
    if (reset) begin
      _T_1187 <= 6'sh0;
    end
    if (reset) begin
      _T_1190 <= 6'sh2;
    end
    if (reset) begin
      _T_1193 <= 6'sh0;
    end
    if (reset) begin
      _T_1196 <= 6'sh2;
    end
    if (reset) begin
      _T_1199 <= 6'sh2;
    end
    if (reset) begin
      _T_1202 <= 6'sh4;
    end
    if (reset) begin
      _T_1262 <= -6'sh4;
    end
    if (reset) begin
      _T_1265 <= -6'sh2;
    end
    if (reset) begin
      _T_1268 <= -6'sh2;
    end
    if (reset) begin
      _T_1271 <= 6'sh0;
    end
    if (reset) begin
      _T_1274 <= -6'sh2;
    end
    if (reset) begin
      _T_1277 <= 6'sh0;
    end
    if (reset) begin
      _T_1280 <= 6'sh0;
    end
    if (reset) begin
      _T_1283 <= 6'sh2;
    end
    if (reset) begin
      _T_1286 <= -6'sh2;
    end
    if (reset) begin
      _T_1289 <= 6'sh0;
    end
    if (reset) begin
      _T_1292 <= 6'sh0;
    end
    if (reset) begin
      _T_1295 <= 6'sh2;
    end
    if (reset) begin
      _T_1298 <= 6'sh0;
    end
    if (reset) begin
      _T_1301 <= 6'sh2;
    end
    if (reset) begin
      _T_1304 <= 6'sh2;
    end
    if (reset) begin
      _T_1307 <= 6'sh4;
    end
    if (reset) begin
      _T_1332 <= -6'sh4;
    end
    if (reset) begin
      _T_1335 <= -6'sh2;
    end
    if (reset) begin
      _T_1338 <= -6'sh2;
    end
    if (reset) begin
      _T_1341 <= 6'sh0;
    end
    if (reset) begin
      _T_1344 <= -6'sh2;
    end
    if (reset) begin
      _T_1347 <= 6'sh0;
    end
    if (reset) begin
      _T_1350 <= 6'sh0;
    end
    if (reset) begin
      _T_1353 <= 6'sh2;
    end
    if (reset) begin
      _T_1356 <= -6'sh2;
    end
    if (reset) begin
      _T_1359 <= 6'sh0;
    end
    if (reset) begin
      _T_1362 <= 6'sh0;
    end
    if (reset) begin
      _T_1365 <= 6'sh2;
    end
    if (reset) begin
      _T_1368 <= 6'sh0;
    end
    if (reset) begin
      _T_1371 <= 6'sh2;
    end
    if (reset) begin
      _T_1374 <= 6'sh2;
    end
    if (reset) begin
      _T_1377 <= 6'sh4;
    end
    if (reset) begin
      _T_1402 <= -6'sh4;
    end
    if (reset) begin
      _T_1405 <= -6'sh2;
    end
    if (reset) begin
      _T_1408 <= -6'sh2;
    end
    if (reset) begin
      _T_1411 <= 6'sh0;
    end
    if (reset) begin
      _T_1414 <= -6'sh2;
    end
    if (reset) begin
      _T_1417 <= 6'sh0;
    end
    if (reset) begin
      _T_1420 <= 6'sh0;
    end
    if (reset) begin
      _T_1423 <= 6'sh2;
    end
    if (reset) begin
      _T_1426 <= -6'sh2;
    end
    if (reset) begin
      _T_1429 <= 6'sh0;
    end
    if (reset) begin
      _T_1432 <= 6'sh0;
    end
    if (reset) begin
      _T_1435 <= 6'sh2;
    end
    if (reset) begin
      _T_1438 <= 6'sh0;
    end
    if (reset) begin
      _T_1441 <= 6'sh2;
    end
    if (reset) begin
      _T_1444 <= 6'sh2;
    end
    if (reset) begin
      _T_1447 <= 6'sh4;
    end
    if (reset) begin
      _T_1472 <= -6'sh4;
    end
    if (reset) begin
      _T_1475 <= -6'sh2;
    end
    if (reset) begin
      _T_1478 <= -6'sh2;
    end
    if (reset) begin
      _T_1481 <= 6'sh0;
    end
    if (reset) begin
      _T_1484 <= -6'sh2;
    end
    if (reset) begin
      _T_1487 <= 6'sh0;
    end
    if (reset) begin
      _T_1490 <= 6'sh0;
    end
    if (reset) begin
      _T_1493 <= 6'sh2;
    end
    if (reset) begin
      _T_1496 <= -6'sh2;
    end
    if (reset) begin
      _T_1499 <= 6'sh0;
    end
    if (reset) begin
      _T_1502 <= 6'sh0;
    end
    if (reset) begin
      _T_1505 <= 6'sh2;
    end
    if (reset) begin
      _T_1508 <= 6'sh0;
    end
    if (reset) begin
      _T_1511 <= 6'sh2;
    end
    if (reset) begin
      _T_1514 <= 6'sh2;
    end
    if (reset) begin
      _T_1517 <= 6'sh4;
    end
    if (reset) begin
      _T_1542 <= -6'sh4;
    end
    if (reset) begin
      _T_1545 <= -6'sh2;
    end
    if (reset) begin
      _T_1548 <= -6'sh2;
    end
    if (reset) begin
      _T_1551 <= 6'sh0;
    end
    if (reset) begin
      _T_1554 <= -6'sh2;
    end
    if (reset) begin
      _T_1557 <= 6'sh0;
    end
    if (reset) begin
      _T_1560 <= 6'sh0;
    end
    if (reset) begin
      _T_1563 <= 6'sh2;
    end
    if (reset) begin
      _T_1566 <= -6'sh2;
    end
    if (reset) begin
      _T_1569 <= 6'sh0;
    end
    if (reset) begin
      _T_1572 <= 6'sh0;
    end
    if (reset) begin
      _T_1575 <= 6'sh2;
    end
    if (reset) begin
      _T_1578 <= 6'sh0;
    end
    if (reset) begin
      _T_1581 <= 6'sh2;
    end
    if (reset) begin
      _T_1584 <= 6'sh2;
    end
    if (reset) begin
      _T_1587 <= 6'sh4;
    end
    if (reset) begin
      _T_1612 <= -6'sh4;
    end
    if (reset) begin
      _T_1615 <= -6'sh2;
    end
    if (reset) begin
      _T_1618 <= -6'sh2;
    end
    if (reset) begin
      _T_1621 <= 6'sh0;
    end
    if (reset) begin
      _T_1624 <= -6'sh2;
    end
    if (reset) begin
      _T_1627 <= 6'sh0;
    end
    if (reset) begin
      _T_1630 <= 6'sh0;
    end
    if (reset) begin
      _T_1633 <= 6'sh2;
    end
    if (reset) begin
      _T_1636 <= -6'sh2;
    end
    if (reset) begin
      _T_1639 <= 6'sh0;
    end
    if (reset) begin
      _T_1642 <= 6'sh0;
    end
    if (reset) begin
      _T_1645 <= 6'sh2;
    end
    if (reset) begin
      _T_1648 <= 6'sh0;
    end
    if (reset) begin
      _T_1651 <= 6'sh2;
    end
    if (reset) begin
      _T_1654 <= 6'sh2;
    end
    if (reset) begin
      _T_1657 <= 6'sh4;
    end
    if (reset) begin
      _T_1682 <= -6'sh4;
    end
    if (reset) begin
      _T_1685 <= -6'sh2;
    end
    if (reset) begin
      _T_1688 <= -6'sh2;
    end
    if (reset) begin
      _T_1691 <= 6'sh0;
    end
    if (reset) begin
      _T_1694 <= -6'sh2;
    end
    if (reset) begin
      _T_1697 <= 6'sh0;
    end
    if (reset) begin
      _T_1700 <= 6'sh0;
    end
    if (reset) begin
      _T_1703 <= 6'sh2;
    end
    if (reset) begin
      _T_1706 <= -6'sh2;
    end
    if (reset) begin
      _T_1709 <= 6'sh0;
    end
    if (reset) begin
      _T_1712 <= 6'sh0;
    end
    if (reset) begin
      _T_1715 <= 6'sh2;
    end
    if (reset) begin
      _T_1718 <= 6'sh0;
    end
    if (reset) begin
      _T_1721 <= 6'sh2;
    end
    if (reset) begin
      _T_1724 <= 6'sh2;
    end
    if (reset) begin
      _T_1727 <= 6'sh4;
    end
    if (reset) begin
      _T_1752 <= -6'sh4;
    end
    if (reset) begin
      _T_1755 <= -6'sh2;
    end
    if (reset) begin
      _T_1758 <= -6'sh2;
    end
    if (reset) begin
      _T_1761 <= 6'sh0;
    end
    if (reset) begin
      _T_1764 <= -6'sh2;
    end
    if (reset) begin
      _T_1767 <= 6'sh0;
    end
    if (reset) begin
      _T_1770 <= 6'sh0;
    end
    if (reset) begin
      _T_1773 <= 6'sh2;
    end
    if (reset) begin
      _T_1776 <= -6'sh2;
    end
    if (reset) begin
      _T_1779 <= 6'sh0;
    end
    if (reset) begin
      _T_1782 <= 6'sh0;
    end
    if (reset) begin
      _T_1785 <= 6'sh2;
    end
    if (reset) begin
      _T_1788 <= 6'sh0;
    end
    if (reset) begin
      _T_1791 <= 6'sh2;
    end
    if (reset) begin
      _T_1794 <= 6'sh2;
    end
    if (reset) begin
      _T_1797 <= 6'sh4;
    end
    if (reset) begin
      _T_1857 <= -6'sh4;
    end
    if (reset) begin
      _T_1860 <= -6'sh2;
    end
    if (reset) begin
      _T_1863 <= -6'sh2;
    end
    if (reset) begin
      _T_1866 <= 6'sh0;
    end
    if (reset) begin
      _T_1869 <= -6'sh2;
    end
    if (reset) begin
      _T_1872 <= 6'sh0;
    end
    if (reset) begin
      _T_1875 <= 6'sh0;
    end
    if (reset) begin
      _T_1878 <= 6'sh2;
    end
    if (reset) begin
      _T_1881 <= -6'sh2;
    end
    if (reset) begin
      _T_1884 <= 6'sh0;
    end
    if (reset) begin
      _T_1887 <= 6'sh0;
    end
    if (reset) begin
      _T_1890 <= 6'sh2;
    end
    if (reset) begin
      _T_1893 <= 6'sh0;
    end
    if (reset) begin
      _T_1896 <= 6'sh2;
    end
    if (reset) begin
      _T_1899 <= 6'sh2;
    end
    if (reset) begin
      _T_1902 <= 6'sh4;
    end
    if (reset) begin
      _T_1927 <= -6'sh4;
    end
    if (reset) begin
      _T_1930 <= -6'sh2;
    end
    if (reset) begin
      _T_1933 <= -6'sh2;
    end
    if (reset) begin
      _T_1936 <= 6'sh0;
    end
    if (reset) begin
      _T_1939 <= -6'sh2;
    end
    if (reset) begin
      _T_1942 <= 6'sh0;
    end
    if (reset) begin
      _T_1945 <= 6'sh0;
    end
    if (reset) begin
      _T_1948 <= 6'sh2;
    end
    if (reset) begin
      _T_1951 <= -6'sh2;
    end
    if (reset) begin
      _T_1954 <= 6'sh0;
    end
    if (reset) begin
      _T_1957 <= 6'sh0;
    end
    if (reset) begin
      _T_1960 <= 6'sh2;
    end
    if (reset) begin
      _T_1963 <= 6'sh0;
    end
    if (reset) begin
      _T_1966 <= 6'sh2;
    end
    if (reset) begin
      _T_1969 <= 6'sh2;
    end
    if (reset) begin
      _T_1972 <= 6'sh4;
    end
    if (reset) begin
      _T_1997 <= -6'sh4;
    end
    if (reset) begin
      _T_2000 <= -6'sh2;
    end
    if (reset) begin
      _T_2003 <= -6'sh2;
    end
    if (reset) begin
      _T_2006 <= 6'sh0;
    end
    if (reset) begin
      _T_2009 <= -6'sh2;
    end
    if (reset) begin
      _T_2012 <= 6'sh0;
    end
    if (reset) begin
      _T_2015 <= 6'sh0;
    end
    if (reset) begin
      _T_2018 <= 6'sh2;
    end
    if (reset) begin
      _T_2021 <= -6'sh2;
    end
    if (reset) begin
      _T_2024 <= 6'sh0;
    end
    if (reset) begin
      _T_2027 <= 6'sh0;
    end
    if (reset) begin
      _T_2030 <= 6'sh2;
    end
    if (reset) begin
      _T_2033 <= 6'sh0;
    end
    if (reset) begin
      _T_2036 <= 6'sh2;
    end
    if (reset) begin
      _T_2039 <= 6'sh2;
    end
    if (reset) begin
      _T_2042 <= 6'sh4;
    end
    if (reset) begin
      _T_2067 <= -6'sh4;
    end
    if (reset) begin
      _T_2070 <= -6'sh2;
    end
    if (reset) begin
      _T_2073 <= -6'sh2;
    end
    if (reset) begin
      _T_2076 <= 6'sh0;
    end
    if (reset) begin
      _T_2079 <= -6'sh2;
    end
    if (reset) begin
      _T_2082 <= 6'sh0;
    end
    if (reset) begin
      _T_2085 <= 6'sh0;
    end
    if (reset) begin
      _T_2088 <= 6'sh2;
    end
    if (reset) begin
      _T_2091 <= -6'sh2;
    end
    if (reset) begin
      _T_2094 <= 6'sh0;
    end
    if (reset) begin
      _T_2097 <= 6'sh0;
    end
    if (reset) begin
      _T_2100 <= 6'sh2;
    end
    if (reset) begin
      _T_2103 <= 6'sh0;
    end
    if (reset) begin
      _T_2106 <= 6'sh2;
    end
    if (reset) begin
      _T_2109 <= 6'sh2;
    end
    if (reset) begin
      _T_2112 <= 6'sh4;
    end
    if (reset) begin
      _T_2137 <= -6'sh4;
    end
    if (reset) begin
      _T_2140 <= -6'sh2;
    end
    if (reset) begin
      _T_2143 <= -6'sh2;
    end
    if (reset) begin
      _T_2146 <= 6'sh0;
    end
    if (reset) begin
      _T_2149 <= -6'sh2;
    end
    if (reset) begin
      _T_2152 <= 6'sh0;
    end
    if (reset) begin
      _T_2155 <= 6'sh0;
    end
    if (reset) begin
      _T_2158 <= 6'sh2;
    end
    if (reset) begin
      _T_2161 <= -6'sh2;
    end
    if (reset) begin
      _T_2164 <= 6'sh0;
    end
    if (reset) begin
      _T_2167 <= 6'sh0;
    end
    if (reset) begin
      _T_2170 <= 6'sh2;
    end
    if (reset) begin
      _T_2173 <= 6'sh0;
    end
    if (reset) begin
      _T_2176 <= 6'sh2;
    end
    if (reset) begin
      _T_2179 <= 6'sh2;
    end
    if (reset) begin
      _T_2182 <= 6'sh4;
    end
    if (reset) begin
      _T_2207 <= -6'sh4;
    end
    if (reset) begin
      _T_2210 <= -6'sh2;
    end
    if (reset) begin
      _T_2213 <= -6'sh2;
    end
    if (reset) begin
      _T_2216 <= 6'sh0;
    end
    if (reset) begin
      _T_2219 <= -6'sh2;
    end
    if (reset) begin
      _T_2222 <= 6'sh0;
    end
    if (reset) begin
      _T_2225 <= 6'sh0;
    end
    if (reset) begin
      _T_2228 <= 6'sh2;
    end
    if (reset) begin
      _T_2231 <= -6'sh2;
    end
    if (reset) begin
      _T_2234 <= 6'sh0;
    end
    if (reset) begin
      _T_2237 <= 6'sh0;
    end
    if (reset) begin
      _T_2240 <= 6'sh2;
    end
    if (reset) begin
      _T_2243 <= 6'sh0;
    end
    if (reset) begin
      _T_2246 <= 6'sh2;
    end
    if (reset) begin
      _T_2249 <= 6'sh2;
    end
    if (reset) begin
      _T_2252 <= 6'sh4;
    end
    if (reset) begin
      _T_2277 <= -6'sh4;
    end
    if (reset) begin
      _T_2280 <= -6'sh2;
    end
    if (reset) begin
      _T_2283 <= -6'sh2;
    end
    if (reset) begin
      _T_2286 <= 6'sh0;
    end
    if (reset) begin
      _T_2289 <= -6'sh2;
    end
    if (reset) begin
      _T_2292 <= 6'sh0;
    end
    if (reset) begin
      _T_2295 <= 6'sh0;
    end
    if (reset) begin
      _T_2298 <= 6'sh2;
    end
    if (reset) begin
      _T_2301 <= -6'sh2;
    end
    if (reset) begin
      _T_2304 <= 6'sh0;
    end
    if (reset) begin
      _T_2307 <= 6'sh0;
    end
    if (reset) begin
      _T_2310 <= 6'sh2;
    end
    if (reset) begin
      _T_2313 <= 6'sh0;
    end
    if (reset) begin
      _T_2316 <= 6'sh2;
    end
    if (reset) begin
      _T_2319 <= 6'sh2;
    end
    if (reset) begin
      _T_2322 <= 6'sh4;
    end
    if (reset) begin
      _T_2347 <= -6'sh4;
    end
    if (reset) begin
      _T_2350 <= -6'sh2;
    end
    if (reset) begin
      _T_2353 <= -6'sh2;
    end
    if (reset) begin
      _T_2356 <= 6'sh0;
    end
    if (reset) begin
      _T_2359 <= -6'sh2;
    end
    if (reset) begin
      _T_2362 <= 6'sh0;
    end
    if (reset) begin
      _T_2365 <= 6'sh0;
    end
    if (reset) begin
      _T_2368 <= 6'sh2;
    end
    if (reset) begin
      _T_2371 <= -6'sh2;
    end
    if (reset) begin
      _T_2374 <= 6'sh0;
    end
    if (reset) begin
      _T_2377 <= 6'sh0;
    end
    if (reset) begin
      _T_2380 <= 6'sh2;
    end
    if (reset) begin
      _T_2383 <= 6'sh0;
    end
    if (reset) begin
      _T_2386 <= 6'sh2;
    end
    if (reset) begin
      _T_2389 <= 6'sh2;
    end
    if (reset) begin
      _T_2392 <= 6'sh4;
    end
  end
endmodule
module LayerParamShifter(
  input         clock,
  input         reset,
  input         io_shift,
  output [15:0] io_actualFeatureCnt,
  output [15:0] io_currentFeatureCnt65536,
  output [15:0] io_currentTotalRound,
  output [15:0] io_currentAccWidth,
  output        io_lastLayer
);
  reg [3:0] currentLayer;
  reg [31:0] _GEN_4;
  reg [15:0] actualFeatureCnts_0;
  reg [31:0] _GEN_8;
  reg [15:0] actualFeatureCnts_1;
  reg [31:0] _GEN_11;
  reg [15:0] featureCnts65536_0;
  reg [31:0] _GEN_15;
  reg [15:0] featureCnts65536_1;
  reg [31:0] _GEN_17;
  reg [15:0] accWidth_0;
  reg [31:0] _GEN_18;
  reg [15:0] accWidth_1;
  reg [31:0] _GEN_19;
  reg [15:0] totalRound_0;
  reg [31:0] _GEN_20;
  reg [15:0] totalRound_1;
  reg [31:0] _GEN_21;
  wire  _T_38;
  wire [3:0] _GEN_0;
  wire  _T_43;
  wire [4:0] _T_45;
  wire [3:0] _T_46;
  wire [3:0] _GEN_1;
  wire [3:0] _GEN_2;
  wire [3:0] _GEN_3;
  wire [15:0] _GEN_5;
  wire [15:0] _GEN_6;
  wire [15:0] _GEN_7;
  wire [15:0] _GEN_9;
  wire [3:0] _GEN_10;
  wire [15:0] _GEN_12;
  wire [15:0] _GEN_13;
  wire [15:0] _GEN_14;
  wire [15:0] _GEN_16;
  assign io_actualFeatureCnt = actualFeatureCnts_0;
  assign io_currentFeatureCnt65536 = featureCnts65536_0;
  assign io_currentTotalRound = totalRound_0;
  assign io_currentAccWidth = accWidth_0;
  assign io_lastLayer = _T_38;
  assign _T_38 = currentLayer == 4'h1;
  assign _GEN_0 = _T_38 ? 4'h0 : currentLayer;
  assign _T_43 = _T_38 == 1'h0;
  assign _T_45 = currentLayer + 4'h1;
  assign _T_46 = _T_45[3:0];
  assign _GEN_1 = _T_43 ? _T_46 : _GEN_0;
  assign _GEN_2 = _T_38 ? 4'h0 : _GEN_1;
  assign _GEN_3 = _T_43 ? _T_46 : _GEN_2;
  assign _GEN_5 = io_shift ? actualFeatureCnts_1 : actualFeatureCnts_0;
  assign _GEN_6 = io_shift ? featureCnts65536_1 : featureCnts65536_0;
  assign _GEN_7 = io_shift ? accWidth_1 : accWidth_0;
  assign _GEN_9 = io_shift ? totalRound_1 : totalRound_0;
  assign _GEN_10 = io_shift ? _GEN_3 : currentLayer;
  assign _GEN_12 = io_shift ? actualFeatureCnts_0 : actualFeatureCnts_1;
  assign _GEN_13 = io_shift ? featureCnts65536_0 : featureCnts65536_1;
  assign _GEN_14 = io_shift ? accWidth_0 : accWidth_1;
  assign _GEN_16 = io_shift ? totalRound_0 : totalRound_1;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_4 = {1{$random}};
  currentLayer = _GEN_4[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_8 = {1{$random}};
  actualFeatureCnts_0 = _GEN_8[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_11 = {1{$random}};
  actualFeatureCnts_1 = _GEN_11[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_15 = {1{$random}};
  featureCnts65536_0 = _GEN_15[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_17 = {1{$random}};
  featureCnts65536_1 = _GEN_17[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_18 = {1{$random}};
  accWidth_0 = _GEN_18[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_19 = {1{$random}};
  accWidth_1 = _GEN_19[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_20 = {1{$random}};
  totalRound_0 = _GEN_20[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_21 = {1{$random}};
  totalRound_1 = _GEN_21[15:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (reset) begin
      currentLayer <= 4'h0;
    end else begin
      if (io_shift) begin
        if (_T_43) begin
          currentLayer <= _T_46;
        end else begin
          if (_T_38) begin
            currentLayer <= 4'h0;
          end else begin
            if (_T_43) begin
              currentLayer <= _T_46;
            end else begin
              if (_T_38) begin
                currentLayer <= 4'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      actualFeatureCnts_0 <= 16'h60;
    end else begin
      if (io_shift) begin
        actualFeatureCnts_0 <= actualFeatureCnts_1;
      end
    end
    if (reset) begin
      actualFeatureCnts_1 <= 16'ha;
    end else begin
      if (io_shift) begin
        actualFeatureCnts_1 <= actualFeatureCnts_0;
      end
    end
    if (reset) begin
      featureCnts65536_0 <= 16'h2aa;
    end else begin
      if (io_shift) begin
        featureCnts65536_0 <= featureCnts65536_1;
      end
    end
    if (reset) begin
      featureCnts65536_1 <= 16'h1555;
    end else begin
      if (io_shift) begin
        featureCnts65536_1 <= featureCnts65536_0;
      end
    end
    if (reset) begin
      accWidth_0 <= 16'h18;
    end else begin
      if (io_shift) begin
        accWidth_0 <= accWidth_1;
      end
    end
    if (reset) begin
      accWidth_1 <= 16'h3;
    end else begin
      if (io_shift) begin
        accWidth_1 <= accWidth_0;
      end
    end
    if (reset) begin
      totalRound_0 <= 16'hc0;
    end else begin
      if (io_shift) begin
        totalRound_0 <= totalRound_1;
      end
    end
    if (reset) begin
      totalRound_1 <= 16'h9;
    end else begin
      if (io_shift) begin
        totalRound_1 <= totalRound_0;
      end
    end
  end
endmodule
module IglooScheduler(
  input          clock,
  input          reset,
  input          io_en,
  input  [7:0]   io_inputOffset,
  input  [7:0]   io_memOffset,
  output         io_finished,
  output [3:0]   io_result,
  input          io_memWen,
  input  [7:0]   io_memWAddr,
  input  [127:0] io_memIn,
  output [15:0]  io_state,
  output [31:0]  io_mean
);
  wire  hw_clock;
  wire  hw_reset;
  wire [127:0] hw_io_input;
  wire  hw_io_inputPush;
  wire  hw_io_inputBufferPush;
  wire  hw_io_inputBufferPop;
  wire  hw_io_inputBufferReset;
  wire [7:0] hw_io_memAddr;
  wire [127:0] hw_io_memOut;
  wire  hw_io_memWen;
  wire [127:0] hw_io_memIn;
  wire [7:0] hw_io_memWAddr;
  wire  hw_io_accEn;
  wire [4:0] hw_io_accSel;
  wire  hw_io_accReset;
  wire  hw_io_maxReset;
  wire  hw_io_maxEn;
  wire [3:0] hw_io_maxOffset;
  wire [15:0] hw_io_featureNumInverse65536;
  wire [15:0] hw_io_actualFeatureNum;
  wire  hw_io_meanReset;
  wire  hw_io_meanUpdate;
  wire  hw_io_meanBufferReset;
  wire [3:0] hw_io_result;
  wire [31:0] hw_io_mean;
  wire [15:0] hw_io_maa;
  wire [15:0] hw_io_mab;
  wire [31:0] hw_io_mam;
  wire [15:0] hw_io_mac;
  reg  inputPushReg;
  reg [31:0] _GEN_14;
  reg  inputBufferPushReg;
  reg [31:0] _GEN_40;
  reg  inputBufferPopReg;
  reg [31:0] _GEN_55;
  reg  inputBufferResetReg;
  reg [31:0] _GEN_102;
  reg  accEnReg;
  reg [31:0] _GEN_103;
  reg  accResetReg;
  reg [31:0] _GEN_104;
  reg  maxEnReg;
  reg [31:0] _GEN_105;
  reg  maxResetReg;
  reg [31:0] _GEN_106;
  reg  meanResetReg;
  reg [31:0] _GEN_107;
  reg  meanUpdateReg;
  reg [31:0] _GEN_108;
  reg  meanBufferResetReg;
  reg [31:0] _GEN_109;
  wire  layerParams_clock;
  wire  layerParams_reset;
  wire  layerParams_io_shift;
  wire [15:0] layerParams_io_actualFeatureCnt;
  wire [15:0] layerParams_io_currentFeatureCnt65536;
  wire [15:0] layerParams_io_currentTotalRound;
  wire [15:0] layerParams_io_currentAccWidth;
  wire  layerParams_io_lastLayer;
  reg [7:0] state;
  reg [31:0] _GEN_110;
  reg [15:0] substate;
  reg [31:0] _GEN_111;
  reg [3:0] maxOffsetReg;
  reg [31:0] _GEN_112;
  reg [7:0] memOffset;
  reg [31:0] _GEN_113;
  wire [15:0] _GEN_13;
  wire [15:0] acc;
  wire  _T_41;
  wire  _T_44;
  wire [7:0] _GEN_0;
  wire  _GEN_1;
  wire  _GEN_2;
  wire  _GEN_3;
  wire  _GEN_4;
  wire [7:0] _GEN_5;
  wire [15:0] _GEN_6;
  wire  _T_52;
  wire [8:0] _T_57;
  wire [7:0] _T_58;
  wire  _GEN_7;
  wire  _GEN_8;
  wire  _GEN_9;
  wire [7:0] _GEN_10;
  wire [7:0] _GEN_11;
  wire [15:0] _GEN_12;
  wire  _T_62;
  wire [16:0] _T_69;
  wire [15:0] _T_70;
  wire  _T_72;
  wire [7:0] _GEN_15;
  wire [7:0] _GEN_16;
  wire [15:0] _GEN_17;
  wire [7:0] _GEN_18;
  wire [15:0] _GEN_19;
  wire [7:0] _GEN_20;
  wire  _T_79;
  wire  _GEN_21;
  wire  _GEN_22;
  wire  _GEN_23;
  wire [15:0] _GEN_24;
  wire [7:0] _GEN_25;
  wire [7:0] _GEN_26;
  wire [15:0] _GEN_27;
  wire  _T_90;
  wire [16:0] _T_98;
  wire [16:0] _T_99;
  wire [15:0] _T_100;
  wire  _T_101;
  wire  _GEN_28;
  wire [16:0] _T_104;
  wire [16:0] _T_105;
  wire [15:0] _T_106;
  wire  _T_107;
  wire  _T_109;
  wire  _T_110;
  wire  _GEN_29;
  wire [16:0] _T_113;
  wire [16:0] _T_114;
  wire [15:0] _T_115;
  wire  _T_116;
  wire [15:0] _GEN_30;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _T_126;
  wire  _T_128;
  wire  _T_129;
  wire  _GEN_33;
  wire [7:0] _GEN_34;
  wire [15:0] _GEN_35;
  wire  _GEN_36;
  wire  _GEN_37;
  wire [3:0] _GEN_38;
  wire  _GEN_39;
  wire  _GEN_41;
  wire  _GEN_42;
  wire [7:0] _GEN_43;
  wire  _GEN_44;
  wire [15:0] _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire [7:0] _GEN_48;
  wire  _GEN_49;
  wire  _GEN_50;
  wire [3:0] _GEN_51;
  wire  _T_138;
  wire  _T_140;
  wire [4:0] _T_147;
  wire [3:0] _T_148;
  wire  _T_156;
  wire  _GEN_52;
  wire [7:0] _GEN_53;
  wire [15:0] _GEN_54;
  wire  _T_161;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  _GEN_58;
  wire  _GEN_59;
  wire [7:0] _GEN_60;
  wire [15:0] _GEN_61;
  wire  _GEN_62;
  wire [7:0] _GEN_63;
  wire [15:0] _GEN_64;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_67;
  wire  _GEN_68;
  wire  _GEN_69;
  wire  _T_170;
  wire  _GEN_70;
  wire  _GEN_71;
  wire [7:0] _GEN_72;
  wire  _GEN_73;
  wire  _GEN_74;
  wire [3:0] _GEN_75;
  wire [15:0] _GEN_76;
  wire  _GEN_77;
  wire [7:0] _GEN_78;
  wire  _GEN_79;
  wire  _GEN_80;
  wire  _GEN_81;
  wire  _GEN_82;
  wire  _GEN_83;
  wire [7:0] _GEN_84;
  wire  _GEN_85;
  wire  _GEN_86;
  wire  _GEN_87;
  wire  _GEN_88;
  wire [7:0] _GEN_89;
  wire [15:0] _GEN_90;
  wire  _GEN_91;
  wire  _GEN_92;
  wire  _GEN_93;
  wire [15:0] _GEN_94;
  wire  _GEN_95;
  wire  _GEN_96;
  wire  _GEN_97;
  wire  _GEN_98;
  wire [3:0] _GEN_99;
  wire  _GEN_100;
  wire  _GEN_101;
  XNORNetInference hw (
    .clock(hw_clock),
    .reset(hw_reset),
    .io_input(hw_io_input),
    .io_inputPush(hw_io_inputPush),
    .io_inputBufferPush(hw_io_inputBufferPush),
    .io_inputBufferPop(hw_io_inputBufferPop),
    .io_inputBufferReset(hw_io_inputBufferReset),
    .io_memAddr(hw_io_memAddr),
    .io_memOut(hw_io_memOut),
    .io_memWen(hw_io_memWen),
    .io_memIn(hw_io_memIn),
    .io_memWAddr(hw_io_memWAddr),
    .io_accEn(hw_io_accEn),
    .io_accSel(hw_io_accSel),
    .io_accReset(hw_io_accReset),
    .io_maxReset(hw_io_maxReset),
    .io_maxEn(hw_io_maxEn),
    .io_maxOffset(hw_io_maxOffset),
    .io_featureNumInverse65536(hw_io_featureNumInverse65536),
    .io_actualFeatureNum(hw_io_actualFeatureNum),
    .io_meanReset(hw_io_meanReset),
    .io_meanUpdate(hw_io_meanUpdate),
    .io_meanBufferReset(hw_io_meanBufferReset),
    .io_result(hw_io_result),
    .io_mean(hw_io_mean),
    .io_maa(hw_io_maa),
    .io_mab(hw_io_mab),
    .io_mam(hw_io_mam),
    .io_mac(hw_io_mac)
  );
  LayerParamShifter layerParams (
    .clock(layerParams_clock),
    .reset(layerParams_reset),
    .io_shift(layerParams_io_shift),
    .io_actualFeatureCnt(layerParams_io_actualFeatureCnt),
    .io_currentFeatureCnt65536(layerParams_io_currentFeatureCnt65536),
    .io_currentTotalRound(layerParams_io_currentTotalRound),
    .io_currentAccWidth(layerParams_io_currentAccWidth),
    .io_lastLayer(layerParams_io_lastLayer)
  );
  assign io_finished = _T_41;
  assign io_result = hw_io_result;
  assign io_state = {{8'd0}, state};
  assign io_mean = hw_io_mean;
  assign hw_clock = clock;
  assign hw_reset = reset;
  assign hw_io_input = hw_io_memOut;
  assign hw_io_inputPush = inputPushReg;
  assign hw_io_inputBufferPush = inputBufferPushReg;
  assign hw_io_inputBufferPop = inputBufferPopReg;
  assign hw_io_inputBufferReset = inputBufferResetReg;
  assign hw_io_memAddr = memOffset;
  assign hw_io_memWen = io_memWen;
  assign hw_io_memIn = io_memIn;
  assign hw_io_memWAddr = io_memWAddr;
  assign hw_io_accEn = accEnReg;
  assign hw_io_accSel = _GEN_94[4:0];
  assign hw_io_accReset = accResetReg;
  assign hw_io_maxReset = maxResetReg;
  assign hw_io_maxEn = maxEnReg;
  assign hw_io_maxOffset = maxOffsetReg;
  assign hw_io_featureNumInverse65536 = layerParams_io_currentFeatureCnt65536;
  assign hw_io_actualFeatureNum = layerParams_io_actualFeatureCnt;
  assign hw_io_meanReset = meanResetReg;
  assign hw_io_meanUpdate = meanUpdateReg;
  assign hw_io_meanBufferReset = meanBufferResetReg;
  assign layerParams_clock = clock;
  assign layerParams_reset = reset;
  assign layerParams_io_shift = _GEN_95;
  assign _GEN_13 = substate % layerParams_io_currentAccWidth;
  assign acc = _GEN_13[15:0];
  assign _T_41 = state == 8'h1;
  assign _T_44 = state == 8'h0;
  assign _GEN_0 = _T_44 ? io_inputOffset : memOffset;
  assign _GEN_1 = _T_44 ? 1'h0 : inputBufferPushReg;
  assign _GEN_2 = _T_44 ? 1'h0 : inputBufferPopReg;
  assign _GEN_3 = _T_44 ? 1'h1 : inputBufferResetReg;
  assign _GEN_4 = _T_44 ? 1'h1 : meanResetReg;
  assign _GEN_5 = _T_44 ? 8'h2 : state;
  assign _GEN_6 = _T_44 ? 16'h0 : substate;
  assign _T_52 = state == 8'h2;
  assign _T_57 = memOffset + 8'h1;
  assign _T_58 = _T_57[7:0];
  assign _GEN_7 = _T_52 ? 1'h0 : _GEN_3;
  assign _GEN_8 = _T_52 ? 1'h1 : inputPushReg;
  assign _GEN_9 = _T_52 ? 1'h0 : _GEN_4;
  assign _GEN_10 = _T_52 ? _T_58 : _GEN_0;
  assign _GEN_11 = _T_52 ? 8'h3 : _GEN_5;
  assign _GEN_12 = _T_52 ? 16'h0 : _GEN_6;
  assign _T_62 = state == 8'h3;
  assign _T_69 = substate + 16'h1;
  assign _T_70 = _T_69[15:0];
  assign _T_72 = substate == 16'h0;
  assign _GEN_15 = _T_72 ? io_memOffset : _GEN_10;
  assign _GEN_16 = _T_72 ? 8'h4 : _GEN_11;
  assign _GEN_17 = _T_72 ? 16'h0 : _GEN_12;
  assign _GEN_18 = _T_62 ? _GEN_15 : _GEN_10;
  assign _GEN_19 = _T_62 ? _GEN_17 : _GEN_12;
  assign _GEN_20 = _T_62 ? _GEN_16 : _GEN_11;
  assign _T_79 = state == 8'h4;
  assign _GEN_21 = _T_79 ? 1'h0 : _GEN_8;
  assign _GEN_22 = _T_79 ? 1'h1 : accEnReg;
  assign _GEN_23 = _T_79 ? 1'h1 : accResetReg;
  assign _GEN_24 = _T_79 ? 16'h0 : acc;
  assign _GEN_25 = _T_79 ? _T_58 : _GEN_18;
  assign _GEN_26 = _T_79 ? 8'h5 : _GEN_20;
  assign _GEN_27 = _T_79 ? 16'h0 : _GEN_19;
  assign _T_90 = state == 8'h5;
  assign _T_98 = layerParams_io_currentAccWidth - 16'h2;
  assign _T_99 = $unsigned(_T_98);
  assign _T_100 = _T_99[15:0];
  assign _T_101 = acc == _T_100;
  assign _GEN_28 = _T_101 ? 1'h1 : _GEN_2;
  assign _T_104 = layerParams_io_currentAccWidth - 16'h1;
  assign _T_105 = $unsigned(_T_104);
  assign _T_106 = _T_105[15:0];
  assign _T_107 = acc == _T_106;
  assign _T_109 = _T_101 == 1'h0;
  assign _T_110 = _T_109 & _T_107;
  assign _GEN_29 = _T_110 ? 1'h0 : _GEN_28;
  assign _T_113 = layerParams_io_currentTotalRound - 16'h1;
  assign _T_114 = $unsigned(_T_113);
  assign _T_115 = _T_114[15:0];
  assign _T_116 = substate < _T_115;
  assign _GEN_30 = _T_116 ? _T_70 : _GEN_27;
  assign _GEN_31 = _T_116 ? 1'h1 : _GEN_22;
  assign _GEN_32 = _T_116 ? 1'h0 : _GEN_1;
  assign _T_126 = substate == _T_115;
  assign _T_128 = _T_116 == 1'h0;
  assign _T_129 = _T_128 & _T_126;
  assign _GEN_33 = _T_129 ? 1'h1 : _GEN_32;
  assign _GEN_34 = _T_129 ? 8'h6 : _GEN_26;
  assign _GEN_35 = _T_129 ? 16'h0 : _GEN_30;
  assign _GEN_36 = _T_129 ? 1'h1 : maxResetReg;
  assign _GEN_37 = _T_129 ? 1'h1 : meanBufferResetReg;
  assign _GEN_38 = _T_129 ? 4'h0 : maxOffsetReg;
  assign _GEN_39 = _T_129 ? 1'h0 : _GEN_31;
  assign _GEN_41 = _T_90 ? 1'h0 : _GEN_23;
  assign _GEN_42 = _T_90 ? 1'h0 : meanUpdateReg;
  assign _GEN_43 = _T_90 ? _T_58 : _GEN_25;
  assign _GEN_44 = _T_90 ? _GEN_29 : _GEN_2;
  assign _GEN_45 = _T_90 ? _GEN_35 : _GEN_27;
  assign _GEN_46 = _T_90 ? _GEN_39 : _GEN_22;
  assign _GEN_47 = _T_90 ? _GEN_33 : _GEN_1;
  assign _GEN_48 = _T_90 ? _GEN_34 : _GEN_26;
  assign _GEN_49 = _T_90 ? _GEN_36 : maxResetReg;
  assign _GEN_50 = _T_90 ? _GEN_37 : meanBufferResetReg;
  assign _GEN_51 = _T_90 ? _GEN_38 : maxOffsetReg;
  assign _T_138 = state == 8'h6;
  assign _T_140 = reset == 1'h0;
  assign _T_147 = maxOffsetReg + 4'h4;
  assign _T_148 = _T_147[3:0];
  assign _T_156 = substate == _T_106;
  assign _GEN_52 = layerParams_io_lastLayer ? 1'h0 : layerParams_io_lastLayer;
  assign _GEN_53 = layerParams_io_lastLayer ? 8'h1 : _GEN_48;
  assign _GEN_54 = layerParams_io_lastLayer ? 16'h0 : _T_70;
  assign _T_161 = layerParams_io_lastLayer == 1'h0;
  assign _GEN_56 = _T_161 ? 1'h1 : _GEN_42;
  assign _GEN_57 = _T_161 ? 1'h0 : _GEN_47;
  assign _GEN_58 = _T_161 ? 1'h1 : _GEN_41;
  assign _GEN_59 = _T_161 ? 1'h1 : _GEN_46;
  assign _GEN_60 = _T_161 ? 8'h5 : _GEN_53;
  assign _GEN_61 = _T_161 ? 16'h0 : _GEN_54;
  assign _GEN_62 = _T_156 ? _GEN_52 : layerParams_io_lastLayer;
  assign _GEN_63 = _T_156 ? _GEN_60 : _GEN_48;
  assign _GEN_64 = _T_156 ? _GEN_61 : _T_70;
  assign _GEN_65 = _T_156 ? _T_161 : 1'h0;
  assign _GEN_66 = _T_156 ? _GEN_56 : _GEN_42;
  assign _GEN_67 = _T_156 ? _GEN_57 : _GEN_47;
  assign _GEN_68 = _T_156 ? _GEN_58 : _GEN_41;
  assign _GEN_69 = _T_156 ? _GEN_59 : _GEN_46;
  assign _T_170 = _T_156 == 1'h0;
  assign _GEN_70 = _T_170 ? 1'h0 : _GEN_68;
  assign _GEN_71 = _T_170 ? 1'h0 : _GEN_69;
  assign _GEN_72 = _T_138 ? _T_58 : _GEN_43;
  assign _GEN_73 = _T_138 ? 1'h0 : _GEN_49;
  assign _GEN_74 = _T_138 ? 1'h0 : _GEN_50;
  assign _GEN_75 = _T_138 ? _T_148 : _GEN_51;
  assign _GEN_76 = _T_138 ? _GEN_64 : _GEN_45;
  assign _GEN_77 = _T_138 ? _GEN_62 : layerParams_io_lastLayer;
  assign _GEN_78 = _T_138 ? _GEN_63 : _GEN_48;
  assign _GEN_79 = _T_138 ? _GEN_65 : 1'h0;
  assign _GEN_80 = _T_138 ? _GEN_66 : _GEN_42;
  assign _GEN_81 = _T_138 ? _GEN_67 : _GEN_47;
  assign _GEN_82 = _T_138 ? _GEN_70 : _GEN_41;
  assign _GEN_83 = _T_138 ? _GEN_71 : _GEN_46;
  assign _GEN_84 = io_en ? _GEN_72 : memOffset;
  assign _GEN_85 = io_en ? _GEN_81 : inputBufferPushReg;
  assign _GEN_86 = io_en ? _GEN_44 : inputBufferPopReg;
  assign _GEN_87 = io_en ? _GEN_7 : inputBufferResetReg;
  assign _GEN_88 = io_en ? _GEN_9 : meanResetReg;
  assign _GEN_89 = io_en ? _GEN_78 : state;
  assign _GEN_90 = io_en ? _GEN_76 : substate;
  assign _GEN_91 = io_en ? _GEN_21 : inputPushReg;
  assign _GEN_92 = io_en ? _GEN_83 : accEnReg;
  assign _GEN_93 = io_en ? _GEN_82 : accResetReg;
  assign _GEN_94 = io_en ? _GEN_24 : acc;
  assign _GEN_95 = io_en ? _GEN_79 : 1'h0;
  assign _GEN_96 = io_en ? _GEN_80 : meanUpdateReg;
  assign _GEN_97 = io_en ? _GEN_73 : maxResetReg;
  assign _GEN_98 = io_en ? _GEN_74 : meanBufferResetReg;
  assign _GEN_99 = io_en ? _GEN_75 : maxOffsetReg;
  assign _GEN_100 = io_en ? _GEN_77 : layerParams_io_lastLayer;
  assign _GEN_101 = io_en & _T_138;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_14 = {1{$random}};
  inputPushReg = _GEN_14[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_40 = {1{$random}};
  inputBufferPushReg = _GEN_40[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_55 = {1{$random}};
  inputBufferPopReg = _GEN_55[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_102 = {1{$random}};
  inputBufferResetReg = _GEN_102[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_103 = {1{$random}};
  accEnReg = _GEN_103[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_104 = {1{$random}};
  accResetReg = _GEN_104[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_105 = {1{$random}};
  maxEnReg = _GEN_105[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_106 = {1{$random}};
  maxResetReg = _GEN_106[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_107 = {1{$random}};
  meanResetReg = _GEN_107[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_108 = {1{$random}};
  meanUpdateReg = _GEN_108[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_109 = {1{$random}};
  meanBufferResetReg = _GEN_109[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_110 = {1{$random}};
  state = _GEN_110[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_111 = {1{$random}};
  substate = _GEN_111[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_112 = {1{$random}};
  maxOffsetReg = _GEN_112[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_113 = {1{$random}};
  memOffset = _GEN_113[7:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (reset) begin
      inputPushReg <= 1'h0;
    end else begin
      if (io_en) begin
        if (_T_79) begin
          inputPushReg <= 1'h0;
        end else begin
          if (_T_52) begin
            inputPushReg <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      inputBufferPushReg <= 1'h0;
    end else begin
      if (io_en) begin
        if (_T_138) begin
          if (_T_156) begin
            if (_T_161) begin
              inputBufferPushReg <= 1'h0;
            end else begin
              if (_T_90) begin
                if (_T_129) begin
                  inputBufferPushReg <= 1'h1;
                end else begin
                  if (_T_116) begin
                    inputBufferPushReg <= 1'h0;
                  end else begin
                    if (_T_44) begin
                      inputBufferPushReg <= 1'h0;
                    end
                  end
                end
              end else begin
                if (_T_44) begin
                  inputBufferPushReg <= 1'h0;
                end
              end
            end
          end else begin
            if (_T_90) begin
              if (_T_129) begin
                inputBufferPushReg <= 1'h1;
              end else begin
                if (_T_116) begin
                  inputBufferPushReg <= 1'h0;
                end else begin
                  if (_T_44) begin
                    inputBufferPushReg <= 1'h0;
                  end
                end
              end
            end else begin
              if (_T_44) begin
                inputBufferPushReg <= 1'h0;
              end
            end
          end
        end else begin
          if (_T_90) begin
            if (_T_129) begin
              inputBufferPushReg <= 1'h1;
            end else begin
              if (_T_116) begin
                inputBufferPushReg <= 1'h0;
              end else begin
                inputBufferPushReg <= _GEN_1;
              end
            end
          end else begin
            inputBufferPushReg <= _GEN_1;
          end
        end
      end
    end
    if (reset) begin
      inputBufferPopReg <= 1'h0;
    end else begin
      if (io_en) begin
        if (_T_90) begin
          if (_T_110) begin
            inputBufferPopReg <= 1'h0;
          end else begin
            if (_T_101) begin
              inputBufferPopReg <= 1'h1;
            end else begin
              if (_T_44) begin
                inputBufferPopReg <= 1'h0;
              end
            end
          end
        end else begin
          if (_T_44) begin
            inputBufferPopReg <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      inputBufferResetReg <= 1'h0;
    end else begin
      if (io_en) begin
        if (_T_52) begin
          inputBufferResetReg <= 1'h0;
        end else begin
          if (_T_44) begin
            inputBufferResetReg <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      accEnReg <= 1'h0;
    end else begin
      if (io_en) begin
        if (_T_138) begin
          if (_T_170) begin
            accEnReg <= 1'h0;
          end else begin
            if (_T_156) begin
              if (_T_161) begin
                accEnReg <= 1'h1;
              end else begin
                if (_T_90) begin
                  if (_T_129) begin
                    accEnReg <= 1'h0;
                  end else begin
                    if (_T_116) begin
                      accEnReg <= 1'h1;
                    end else begin
                      if (_T_79) begin
                        accEnReg <= 1'h1;
                      end
                    end
                  end
                end else begin
                  if (_T_79) begin
                    accEnReg <= 1'h1;
                  end
                end
              end
            end else begin
              if (_T_90) begin
                if (_T_129) begin
                  accEnReg <= 1'h0;
                end else begin
                  if (_T_116) begin
                    accEnReg <= 1'h1;
                  end else begin
                    if (_T_79) begin
                      accEnReg <= 1'h1;
                    end
                  end
                end
              end else begin
                if (_T_79) begin
                  accEnReg <= 1'h1;
                end
              end
            end
          end
        end else begin
          if (_T_90) begin
            if (_T_129) begin
              accEnReg <= 1'h0;
            end else begin
              if (_T_116) begin
                accEnReg <= 1'h1;
              end else begin
                accEnReg <= _GEN_22;
              end
            end
          end else begin
            accEnReg <= _GEN_22;
          end
        end
      end
    end
    if (reset) begin
      accResetReg <= 1'h0;
    end else begin
      if (io_en) begin
        if (_T_138) begin
          if (_T_170) begin
            accResetReg <= 1'h0;
          end else begin
            if (_T_156) begin
              if (_T_161) begin
                accResetReg <= 1'h1;
              end else begin
                if (_T_90) begin
                  accResetReg <= 1'h0;
                end else begin
                  if (_T_79) begin
                    accResetReg <= 1'h1;
                  end
                end
              end
            end else begin
              if (_T_90) begin
                accResetReg <= 1'h0;
              end else begin
                if (_T_79) begin
                  accResetReg <= 1'h1;
                end
              end
            end
          end
        end else begin
          if (_T_90) begin
            accResetReg <= 1'h0;
          end else begin
            if (_T_79) begin
              accResetReg <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      maxEnReg <= 1'h0;
    end else begin
      if (io_en) begin
        if (_T_138) begin
          if (_T_156) begin
            if (layerParams_io_lastLayer) begin
              maxEnReg <= 1'h0;
            end else begin
              maxEnReg <= layerParams_io_lastLayer;
            end
          end else begin
            maxEnReg <= layerParams_io_lastLayer;
          end
        end else begin
          maxEnReg <= layerParams_io_lastLayer;
        end
      end else begin
        maxEnReg <= layerParams_io_lastLayer;
      end
    end
    if (reset) begin
      maxResetReg <= 1'h0;
    end else begin
      if (io_en) begin
        if (_T_138) begin
          maxResetReg <= 1'h0;
        end else begin
          if (_T_90) begin
            if (_T_129) begin
              maxResetReg <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      meanResetReg <= 1'h0;
    end else begin
      if (io_en) begin
        if (_T_52) begin
          meanResetReg <= 1'h0;
        end else begin
          if (_T_44) begin
            meanResetReg <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      meanUpdateReg <= 1'h0;
    end else begin
      if (io_en) begin
        if (_T_138) begin
          if (_T_156) begin
            if (_T_161) begin
              meanUpdateReg <= 1'h1;
            end else begin
              if (_T_90) begin
                meanUpdateReg <= 1'h0;
              end
            end
          end else begin
            if (_T_90) begin
              meanUpdateReg <= 1'h0;
            end
          end
        end else begin
          if (_T_90) begin
            meanUpdateReg <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      meanBufferResetReg <= 1'h0;
    end else begin
      if (io_en) begin
        if (_T_138) begin
          meanBufferResetReg <= 1'h0;
        end else begin
          if (_T_90) begin
            if (_T_129) begin
              meanBufferResetReg <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 8'h0;
    end else begin
      if (io_en) begin
        if (_T_138) begin
          if (_T_156) begin
            if (_T_161) begin
              state <= 8'h5;
            end else begin
              if (layerParams_io_lastLayer) begin
                state <= 8'h1;
              end else begin
                if (_T_90) begin
                  if (_T_129) begin
                    state <= 8'h6;
                  end else begin
                    if (_T_79) begin
                      state <= 8'h5;
                    end else begin
                      if (_T_62) begin
                        if (_T_72) begin
                          state <= 8'h4;
                        end else begin
                          if (_T_52) begin
                            state <= 8'h3;
                          end else begin
                            if (_T_44) begin
                              state <= 8'h2;
                            end
                          end
                        end
                      end else begin
                        if (_T_52) begin
                          state <= 8'h3;
                        end else begin
                          if (_T_44) begin
                            state <= 8'h2;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if (_T_79) begin
                    state <= 8'h5;
                  end else begin
                    if (_T_62) begin
                      if (_T_72) begin
                        state <= 8'h4;
                      end else begin
                        if (_T_52) begin
                          state <= 8'h3;
                        end else begin
                          if (_T_44) begin
                            state <= 8'h2;
                          end
                        end
                      end
                    end else begin
                      if (_T_52) begin
                        state <= 8'h3;
                      end else begin
                        if (_T_44) begin
                          state <= 8'h2;
                        end
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_90) begin
              if (_T_129) begin
                state <= 8'h6;
              end else begin
                if (_T_79) begin
                  state <= 8'h5;
                end else begin
                  if (_T_62) begin
                    if (_T_72) begin
                      state <= 8'h4;
                    end else begin
                      state <= _GEN_11;
                    end
                  end else begin
                    state <= _GEN_11;
                  end
                end
              end
            end else begin
              if (_T_79) begin
                state <= 8'h5;
              end else begin
                if (_T_62) begin
                  if (_T_72) begin
                    state <= 8'h4;
                  end else begin
                    state <= _GEN_11;
                  end
                end else begin
                  state <= _GEN_11;
                end
              end
            end
          end
        end else begin
          if (_T_90) begin
            if (_T_129) begin
              state <= 8'h6;
            end else begin
              state <= _GEN_26;
            end
          end else begin
            state <= _GEN_26;
          end
        end
      end
    end
    if (reset) begin
      substate <= 16'h0;
    end else begin
      if (io_en) begin
        if (_T_138) begin
          if (_T_156) begin
            if (_T_161) begin
              substate <= 16'h0;
            end else begin
              if (layerParams_io_lastLayer) begin
                substate <= 16'h0;
              end else begin
                substate <= _T_70;
              end
            end
          end else begin
            substate <= _T_70;
          end
        end else begin
          if (_T_90) begin
            if (_T_129) begin
              substate <= 16'h0;
            end else begin
              if (_T_116) begin
                substate <= _T_70;
              end else begin
                if (_T_79) begin
                  substate <= 16'h0;
                end else begin
                  if (_T_62) begin
                    if (_T_72) begin
                      substate <= 16'h0;
                    end else begin
                      if (_T_52) begin
                        substate <= 16'h0;
                      end else begin
                        if (_T_44) begin
                          substate <= 16'h0;
                        end
                      end
                    end
                  end else begin
                    if (_T_52) begin
                      substate <= 16'h0;
                    end else begin
                      if (_T_44) begin
                        substate <= 16'h0;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_79) begin
              substate <= 16'h0;
            end else begin
              if (_T_62) begin
                if (_T_72) begin
                  substate <= 16'h0;
                end else begin
                  if (_T_52) begin
                    substate <= 16'h0;
                  end else begin
                    if (_T_44) begin
                      substate <= 16'h0;
                    end
                  end
                end
              end else begin
                if (_T_52) begin
                  substate <= 16'h0;
                end else begin
                  if (_T_44) begin
                    substate <= 16'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_en) begin
      if (_T_138) begin
        maxOffsetReg <= _T_148;
      end else begin
        if (_T_90) begin
          if (_T_129) begin
            maxOffsetReg <= 4'h0;
          end
        end
      end
    end
    if (io_en) begin
      if (_T_138) begin
        memOffset <= _T_58;
      end else begin
        if (_T_90) begin
          memOffset <= _T_58;
        end else begin
          if (_T_79) begin
            memOffset <= _T_58;
          end else begin
            if (_T_62) begin
              if (_T_72) begin
                memOffset <= io_memOffset;
              end else begin
                if (_T_52) begin
                  memOffset <= _T_58;
                end else begin
                  if (_T_44) begin
                    memOffset <= io_inputOffset;
                  end
                end
              end
            end else begin
              if (_T_52) begin
                memOffset <= _T_58;
              end else begin
                if (_T_44) begin
                  memOffset <= io_inputOffset;
                end
              end
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_140) begin
          $fwrite(32'h80000002,"bn abmc: %d %d %d %d\n",hw_io_maa,hw_io_mab,hw_io_mam,hw_io_mac);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
